XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ZJ]?��oP�ön����l�b�;�}�o�'�n��߭a��ƑD��p�	Goƪ�Sb)-k����N��l�	S���m�t�Q�t��G������hlU�JQ��:f�������'ݼL���E��W� ��怸���%	�:u���Ea��L�.��j8	5d�r�HLg� r���E
�"��3��'��;��Q!�z�c{h.]Q�y��Zoh�z�9ͬ�,�d��>5)^��V~%ʎR�'(���Z���V�]��z����t	���\$�k��tt4Q��IN��C���Rҏ� GյZ����	5S� 8�M���vm��6���������2�:����O>��HX�<�M�8��}҉��&�À1��&.J�^[����H���rZ��ԧ����0>vƵ�[Y�+�V,^:��g9g+x�����G_�q��o���"�H�O��y��C� ��tEk��S���ɤ���yIR�Ǒ<nL/7	{MH�Q��L�Jr���*�mҁ����Nc��t�A�v�+�O*)�ȓr?NH4v�D\�e:��})q�����X/]E�+(�[�-�]��R~�1�ש2*�y@]=ʸg��vM�&�*D+T�`��z��A�eC�R�k���\�l�с%��57��Bw�Z��+p�k�R'�=b���49g��l��1�E�@�(���h���J4z-]�bK�:�����(��&��zz�n�Π���A<IKU��>�J#\�ҵ|��aS>XlxVHYEB     b88     3c0!:u`�>�yI��l$��@��k�����o��7$�8��ғ4�í��G��r�A���
CW��5j�mݽ�'|Sa<���N�v���8cne;���p�$�c;��%�ܝŕc�7��sg�?�#�*�om�FfhvRh��M�SU�1)��s�
? sP� �Q�VY�I>
M�*�2.:���ɒ��)(Ut�F�8�4fW:��[-��๡���0u���H�l����
��@�&���M]
����0����s��dH��"K�,�ICG��g֪�sI�0�~�COd�*��F�  ��"��j�� g��<���.	;e�����҇
��H�7?4۰n�0�-R*�^�� VEK�KnO���f�A�T�j���D�i���6>ڃZb�wi�����)` ��T��-@��:�����3C0H��ǜ�NKzym�:��Sę�@�}#d�<��Lu�>�Y���tI*H@L�R/�!B3���̙<9�>�;�]��v��pה������6	���{=9���F�����	rcU �9�;G��A`\�&�dU����/��I�VX�"�7�;��
J��˲ x����3a3�|}�gLz%ئ��������-yO�1��:���W�<���ٓy6`�E3�Z�@��`T�lwiќ���~�3���'G�n��S��̳ӏ��_��T{�K����/�`���WkTx�--$�@2V��/��!�r(��ْx]��_L�9~"S!)�V
w�� �O�����ꔽD[�y��#��X�:����d V��V���Ϛ��ݶ�nӣ�J��
(��@�S�\q���*�֜���	�E��2��½xáo�ϭ��WXd+BUrzl ����J�37�p��v�ӗ$y����aD����~����'d�;U�/��W.�$�yψgh7<"E�`��Cy;M�1�<����o��V�3I�R�T��