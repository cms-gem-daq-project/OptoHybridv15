XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)U��	�K&n�/�V�k"�)k�>y^�P���B��r*��Ԯ5�v��rS8[����;��|��A����M��d�(W� �&�
)b`�	�8^&;4ZdiB���X�u=��RY;\�)	#���咃�|]���RȒ��sz��a�1aG�6�'�>P>f��E����t\��G�S�C�r���+Rp�׃���ľ*Ŷ2�Y*�����寖o��i7��8���a{
��C�w2�q��w>*<�*�Of���T�����	lF�96�I���Ǵ
�"���Y�L����K@,��8X8� N�$s�p0}���Z�1����q����gj`�y[VŚE�m0��>!�E�F�I$p�00 m�|y���4_�4��b%e���e��|ꨬ��/�,�}�3��4�C|�#,%�<�MA�gȡ�e�ۺ���ϋ�Ѥ���C��C����I���{^��C�XBV�i$dj��/�4I���V���x,���6���%Nj��K<�JrS-��8z�2�/���j��APɩ��w��X�wc�] (��խ�s)(ۑ�D�1�8K�R
�
O�[�}��m=m��h?^����?@�ۃ����:#�ݻ���6L���]��F�c�U5$���z��;��U�f7����(�یQ��2�a��♟�]�Q���8v׋�%Z��l@f^`$�O�./A���m���}��{�5����v=c�.�a��Q�`���P�~_q�f<��.�(������b)IXlxVHYEB    3c92     900�]%���W��0�wd+N��-���,>Z��+l��h�Z��2E:C��ww��z~��pf9���xkX�ip���|ơ�vD	M�p=r���>�U�7F�o��V��Ng<ۖ���6��+v3���J(�΂E��,��Ĳ[��Ǟ�����]&�f�!�w�}���r��X��k��iL�1$��4tA��^�͝6��8�+��v{�o�f����ӷ�{������l:-���@˱�R��Rw*|���ܤ���^��G�+)g��,%�^e�Z���\�:�P�?��H'ú^8���B���XI�3��q��7�¤y}	��ȏ�$/��{���.����G�o�2/u��kb�l��!6�9AR����
��7'�xu���: �ۆ>�x��bh��O�Ō���J����*��!K��1.��C��<lӸ;� W|t��g�AF��c^�|J�ا�y��ՍI\C�MG�NX���Q������b~��C]�Cb��8�ĝ&=��]��e��CM�:kl��İo���N��*�{�}�ʛ,: V8I��p�\B4���!�t����=���(Zt�.��.L�����#�Z<-�8��Pn�4ʃ]]I(���zJ|ĘM`t�{
�*\��}y�[�d���@��j���vP��z/�7��Ҩ��]n�;���ʑ,��76�ث���|Y�N9bgv�xʯ@�l'Q�6��[�]_���ag��%�?Qp�j���3m T`���8a�-�$/4��I?nC:ޝ��@���a�%��E�5&!s�G��r��k8�1	#�Pät�����ۼ�z~�#r�J��
x�_�`X�[T����-6���V��q�g<a�!��d��M6�X�m ��>x:�)a�wY��,)�F��2�Ɣm@��|�@��qK�Bl���~li4s�^�㨗�%y�ݤ����b��^����݀��8�����>�Ǟu!�<r���ȼ��ǳ�QI	��^u���݋F	�y aZ8��*� �fOp=��a��s�����ܦ+ FR��i��>�c^m��%�qCyn���k���Ţ�e��gqH�o ��̨g������sT��G����.�l�|E��l�[�C���WF�A��1��vq�qC�w�ic����ɸ{"E	f��w#+�8��6�3-��d
M�%�7/�|�^S���[VY;)
27�@���ܒ:��O}���C��[�؀2b��N,d�@��p ��ʅ�I��Q���ו�n#t11�3��9h���$�w������h�e��T9�#��'n�6��9@�l�J�Ē�fĐ-�w�b�mʩ��j�'���y!���=[��BLx�`�?��gt2�����р�o>xh���)�QX��&�30��V�M�H%F�g���*�oP�,a'�tm�d�K6��~ov9)<��ު�h�X�!�K�:-jޫP.�X��(�>��N�}<��\�YPQ%-�����t'�V��K����i�r^�����(����L�u��u$ �r����ˀa#�cT����)ʦ7�E��o�K�R,Jvt�J&��v��Z��ZCk�2u���kTz�m���p	@��a��%��y��B�V�D�x�3�t_�=GW�(Hׄ����e�ٜ�GH�Gkc��v��~Ǫ�8w{!��C ����$A��E��P.ڴ�����3�&�ۡ�%9��� ���E��r��	ŕ���Ge�/w�	�"(#k���5��5�j\��uy�f�p�RI��M�:N7x�ׇ˼)��a3ڱ8d?� �ƶ���	`P�yz���B���2��*U]���ww�k��T��|.�E��=�2r�$x ��EQ@�b��Xt&!��� 2����,ٙR�ހ{�﬿���@�X:���=���/�k��|_���UD+����/� �| ���\�֢Vi����=�j���,	� �d�S6[�l���nٹ����D,��	鯺K�
�lz4���Jl+=��A�G���[�WL�i3&t\�&,KΙ�L�����X4��`��8)�:�q*�j�e��c�ϖi��k��PZ���c���~��OK�P}�v��_�p��C�I�O�Ա?��Ac��y����Vd�<:�乫�MQ.)�*)�8c�盻N�P�*2�2J�K�7�"7�kS�Ĉ`���B�A�b��:��m����.ш�¸?�Th���1��>	g1��l!|>xv�h�9�JH�RO|�<Ԕ�o�c