XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����MMGu��Ҽ�&/�+���N|������<W����z�$Am=,�V�?���r#�Kמ���v�s�tJ�H�Z���xw��Y?sd�	���<X,<��x{?��ե���d��C�4���n���`�+'*����o�/�`�i���8�a��@�î$�4H!�q�狦r�C�N�B�u*�>}]M/���!��߬w��Fx4*�VEZ�%_sf'�(�>�\��y����	"(�Q�0��_D�-�'j+��K�غ ��OYE=�	OL��)TMt�`_�7�L�â�� !VԸ5�"OR�������Mj~+�E��K$M5�W��#*H������A^��&dɕ�y�.�D<}�P����.m�|�)%`7*�p��No\���F��F�s�6�@+���Y_�e��BƟ�_�
��ot"���rL�d�i��c��:U=��eu��a@d�/L�+�k�\jS���v�0pB>���v�W����;EW�`����pf�kFChl�۬�Tlw�Z���a�i2��g�e@��U�U�۬i�S��A������^��k�z�����Hג��a��UbH���1ɐ�w����	�<���F�r���6.e�&ӡu�/�D�䨩|��@)��zxN,%��!d��v,H�0y���.�̘A�{�9^�kR���eh�_S�}ͅӯ.ض���Te� ���L��Ԫ%vV���IM�6��%�ܮ���zgB�G��Cve>NH�;ld�.D��]�-�`yl����XlxVHYEB     b8b     3b0����p��ZҊ��ߒ����g2 c���Ye�8h����юY/�[<{6���xXP]h�G2����O	�ݫK����VˊeB���G�הR?baA��˯��N���P�;V�veP�ۚs�*kUs���2�;��뵽�m�x 4�uv�X���Y��/E�]�D�qx�A���'p*.�r���6$ҬW�0{W�� ��j =3���_����x�8w�9�g�\,�֔ͱSu߲�Z�txɎw�Kʇ�p��<�� j�M�6�U4X�YnGfpގ}r�yc
��6tbr5��a�S/��Q�'�-��z��_6Fgp��H����v�n����6�sc����z{�o��Y�x���r�+,]�����G��G�d"����,�6�s��|f����r8<:W�����δixF
LX��Qh����@�J���_�BQ20R7��֋��S9+#�D]凋�]�W8�P�=7����ݽo:;�^�ߋ=���Ls8�qC�>�;���^�K�HϦt��7#_��uDTҖ�~C���X�y�������
�wN/z�T�xȢZ� I�hjh%֪���o��kY�4���pJ�mj����m���W2	��beF�Z�h�Ց�[�D��P�@xWb4���>Is׬������e\�oelWM�AAȲӃ_O�a��V���&�{�p��y��w�)W_�)�d���˥��]�]v�����	v,��3��r�u���t"q ��1Oy�U^�ԗ��]Tt֋ �*?��P�"�~G8���XO������W�J�/04Bg;��`��]��v�o^=%��6R�Ƣ������lP���F ��r���%��)����bV:�@4�tu�Mi#F����[�/aM�:r�!9�%*��)7h�K�?�?�q	�ƶY �tn��^�-��n
�D� �03�{�^�-