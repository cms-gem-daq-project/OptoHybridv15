XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&z�d����-���{�:�lj�z�
�6��N#��7e�6M�E9]��g `�}?p9G��ڴ=5R�-[�!������(�����L�L�9��mQ�x=��b����x�B�+��#V�&\������D������|�� ��6WP �8������ 4Բ�k�S�(�(���j� �Ts\z�p0�0�V��>W|w�klE�QE �_�>��գ�[~��K��zK��J��I������&i����d�%]pD��ȣ���&���և~�>�1�	]�0:�:�z�lfۇB8�I�,��w�ـB�o�> Og�Ӯ��Ͷ���L���an��Ln�)ncj��u��e��2���ձ����:��W7G�ZA�R���4�BpᩀF�m,fP�ꯑ�ƾZʉfa�$;����hA���6#�9���������еM<�G��/ʣ%�N緾�y[�-\��>�a�|6v��`u�f!`�z��^�[��^Վ�n���!��i�:%�D͍�5=��Mm3!�[r���h���*!Z���jw�J��i�-�tTD��ZQD�O���xh�XNs��eT�y��	�$?Ck�M����X�lH6�Q�����V����t�^�7FDo<n�2���u�,`k���m-�E?�Y�У.Ɠ' x�WS uS6����|
Ů�rO8ڏ�S�HX��������SK�0lO��Qjm���;��k�R�j)����U� �"���9<����
,�w~����XlxVHYEB    1621     410x��c����d��}�����9N�Z�*�!��C�K˷O��OU$����lY[\5n?�d0�5!�[�}���[G("�
c
�܊?4�#pX� �¼��A�lM&?�K�1��%+���K���!�\�:��6��b�e���r��Wh�;�_���v�������gUSW�\��ӏz�z�КַL-�B&�:���w���'��mJ�m1�:뿌'M׺q�rz,�C�G��%�}<�]��%�֯�PL���7i���Jw�]]�،�9.��Iz�1LPw|`��7%���S֫6)��"C��̠�{�k]��-��DOJ΀+��i��y�+�xr��t��#��Q�e�Dڠ�1C�zZsWmt0a�'?�ʝ�͐=0���dbR�������!ɗ&,��e�@�n��3��M�ge �]�!&Xk��%�@��0��w�O�2�;���U�`ŬZ��Hdv���p?��}�wJZ(	�C��$��4x�^�9��j�/���B}��$��՘Jo�} %��F�@c�/��V�uZN�/ t���R��sc�"�Uvq����܅5�6ȫ�'uɬ���3�Kc]p�4����a#5��T���hA�3�E:q7�ص���&ፒ����.�#��p#��YA�d�F":\%O5�Ntce�[�<.��b1"_mWt��AiAO"z��OOE8q��.�9,���ǯ�TߘO��s��Y�Q��}ۢ��=��g;�v.Cg*��;~msu��U�Ű�D�0�����b���� ��Gϻ"��g����7�\�5G{ju��5�V����Ȇ�g5ufH��j�7`}�
��a����5�Tl��fP6<"VU%��%���/�����g��CU�x����GL�����伎�|�%�@�	G��I=�y�cM�2)��w�sқzԆ�MF���X�����&x�ޞ�n�Ҏۑ�����>d���b�"��3E�y���

܈s$
$�Sz+|xp+)2c6��f6��
�țc�