XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�Wd ��*��rp���KD1�:�)�u��O�F�2��Wb�I.ֺ���#R�@?����.&h#��:�Ȳ:}r	�0_�YR{�M �~<ُ�!���X�ls��}��?�89��B"TqH+�$֯c�Ʀh���,πT>C��7(@΃����D�c�1�s����@j�k
�n{�'�t;"6̷������y��+���n��>��%ة�,��)�V�%���6��Z�s�d�`���_/e�u���70/	]���	�,�+��U
��34��,1D�75��D�F�B&ǐT��{�mVO�Pw���a�6Q�
��h��n�$�Ͽ������3�*SR G�;8|�S��6��:��o�t@��s�9,=�� }x�o�V#��9A�'˳%a� ��B�7�Z�RS�XR͜�?v��m#��5:���/|y�D4����_<����>m�qx�c��T������9�@�N�K�+v^Q�y�6tE��gYɊ��~	UM��NT"H=�:@Q ��3�A��z��y�t���uT���3hi�L�6mR�А�d���Y��]$9��Ģ3u	+n��~�>m��F{x]��)�v�	��0�|s���z�GC�7�����Z�� �#MBš�J��;?�P��JUFJ��f��R��t���JiQ>�\�U�0Bo����<7oN�/�Thj˾#FQ��j�L/%<3>�Qa�)�l���D^��h��1̚���{����N'�YB��"� ���}Q��B:��ͪv:�C�Sn XlxVHYEB    166e     400]�Z�K!�`��Mn����*��Z�a{CS=�س��·\�:÷�Z�w����'i�6jlt���Py�2;��JVN~5c���G�ݔ欅I��J����#a�؍O[I��#hjf�^>��JC3S��_ ���JN�8�/8zd�L����Eq����s>���������{������,^\��~~�=MF�G��f<�8As��\qt�U~!��Ձ��-��QuPN��{�!%7�.��[�|���p�&/i��:��9��y,���Ns�G�,S�iu���[_��\ƞ܏G`.֢���}����N������'T��|��J��Ǩ׽h�_�e|:����r�A�Ŕ�iV.JU�l����W�CYB^K�	�_y�ۢli�ԧP��:��4�,�p��Ӧ��-�&e��9}�~������DJ�[v��>�~�t�.���K�-�)��[*N3_g�/r�װ��b�~L�T��zd�5�J�� ���N�'� �����9��c���&}����w��D�����߱���ћ����ꡢ݀ծy�l��C����[��%*���j���<`l �Qg��U/nʶy
�_S�"�tNP
;j>��>��]����~��"���5g:z"v�CQ�DbX5c�C]7d���٧G��Xl�e3�3�'jK�����ҒZ���Hb��S�:��d3h7=&�	D�����(��� �����E��븫{���f`��8��ٰ�H�Nۂ{��
����>�`I�a�q6|�����2�I٬�*z�/�%6����X��5n�͘��g�v�3OK�ֲ���o��#�|ً�8�2�`�8��1���Oq�ǂ�*")cb���'Pw/�*(닎�%Ϻ4���Կ�m�M��j��$��>��� ����%־�����GG-ti���~D#�Y![�������+Mt.$o��2���xҝ�N�Պ������{�ۘ��VE樑
�'E�gm�U�Æn��/��^ʆ��`ڏ����brp╷��