XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�M��WQ��b�7�h�m-#�ϣ�Ujܬ�3�<�yl��@I:�!�PB�����a|Y^J_v\8�0����u�0�g6 vj']j>����v�e]���2����`�f}�KV:JJe��x�UPK!}ƌ4�4���%�SH���˅�����˓��/[������7��.f7vK��(�,��UU ��[���I�gNqҨ3�*���M�F�B�ݏԻ�h�LW�.���� 3�����J-�Ԥ��M�z֎�c&�����q�7����U�*ߖH��}��ߚ���[�.��~��
W�*��6�&�<��0ݑ?,�]s�R):#�CC��܊Z� �p�f[�¾�R���Ơ�]�{fDX��egO,�dĘ�I��꽀'�����σ�"D
7:���7"���G����!ym|a"u8��0��>i&#�h+�[ˎ��/���R2�IC2$<���`)[�9���.�0���S�V�"P��(���AY�E���J���1��H���ŜQ�J��I����<6�L�A�(���'���(ߡ�R��o:U�Ѳ��aL���
��n�~K�Y����6�����RA�q���I��ʷ��;����$�u=�|�>�,�[�%�<ȯ���mX��ka��>P�݊`�� �٫+�W��t)]u8��rg�-(�Z�
_��k�~JB6������c�/u�CD�m~����F�~ؠO	��aY`_���-�o���������d���/�������=�j跛�XlxVHYEB    11e4     520�Y�u9�L{�2~Uj�Q]s�t����I��bEg��&s�����]����i1h��Ox�դ��|�U��MR3� �ݗ���Lj�e�s�=`}�I�����ud�ܣ���-B�*�� �F��Mc3��xGhO�Rx�y��涐���Q�������'��"���3]uk���&�'
Ͻz���5���	�/���t�v%�"��;u�w��E̢�������S�F�������+w`A�.7��]��!�~���G�b���r�P4�s�A	��R���OU�*�}?�6�R��Mˇ0,��`;�
 �Өʀ,����ș��Y�"gz�����<p/�U2C�����qk�@C�H���9����q9/�ԗ�kn��8^L��½<���t�>�0b��.O�8H��&������h���Y8�#�
�ԟF�d��m���~4�b3Y����N���"��[�S��%��6�Dw��ئ�4ӳhQc��@bh��`o���ߕ�Z@@�B�R�Wz��������S�c3*�d�� ��6�z�D�MP?G����zc��$�N�3(�z���e|���B\�Lѕ��թ-��t�ƛ���ً��6�e�	ې�J��Y�R�C�j�{N�D��껾���Ts��@��Q�zG��V+Ҷ?��L���v���rI�3�V��xJ�(�p�醖~�h�d%g|���/D��`)���d$l��|y�'u�J:��|���U, �;��~2��{��_˕Y�6�5��.�0VCo2�� }��l甖�u��b�Q`n�7;%]���}ڶ��^�e<!TE��D�{�-{��d����]���
�����&p�����U��!f�%b����紐p��t�T{"�\�M���끃��[����M��a���������t}�$p ���^����M�R�k��=`�-��[�i�*%b���m�B�Q�T��.K��s���w���VŎ.�$��B�B
��%S�s�=�4����H�H�����\�c���ך���L��|�Y_�]���$͋�2�Ŋ��>����c{�R��p��e�� E��o�l*|�؟�:Al�Gz�?=W.�6P�Tũր��/��6=%)�/�`$�_�S_4�(%d�9Dyٛ��2�`�E�"�oZ�n _�(�7��cvᅏ*�^o[�����+�S@U.gv�lE9m�:33r�O򋿮��R�1��~�I�5��Q��S�)j߾>�z�� gq�?.�j�+�.��w5F���X5����N��x���b����vX�L�