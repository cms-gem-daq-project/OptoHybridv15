XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}J��v�*a�!E`��4-�^|�U��'Ի�|��3=�X� G�Xi��	���SA��G��*�Jx)��&����wK��ߴ"�J/����V�Q�M�w���IC ���q0 ���K�]X��5���>����I� ?��m���NbU�8��3�>��u`]�ڗ����4i$6��RDpO�q�^�����IJhy�e�:討i�U�1�҃�{���I]x�v�����?JyQs� �Z4����#�N��m�f�ɲ3v}��wm�%~�O&���%���9�[�Ur�;��|���~s? �E�P#�-�0�VJW��1�2QV'th]�&��ȫ�7��BW�D�Wqٶ0܆#�����I�m�9��x�x76'��z�zM�
[�q�<�e�;8�[�'�XY����j��Yp��`ر�
ok��G3fi~�
����P����D��T�iQ�Iq�"sޛ��JpgX?��wI�����Ch���P��7��\�յŹ�ª(�ɽO���C���0e�H庚�S��bm�4����gj���ߠ7_�Ք�ۧ��^�.�'_��S���ߋ��i����C,�� d*�^�e](M���jE�۾�^��
5�,=lR !kݣF�Ex�l�}�02� a�]��G�Y���������О������SWt��)� -�&�������.L���
�
����(�6j�˧i�	{g��h�e�����(�ˢK)Z��ۿ�
m������H'\�lT��;ʃШ�\����QT�Јr<XlxVHYEB    9b67     f50�8W��28UM�����P��G�*7i���R��/����Â�v�o\RG�Pv��>�	Ç_8o�y���5?���t۹���6�>����_k;9W�寓W>���(��gI=�Z��4`E.]p���jt�e[f{��J�.����p4ß��UgQ��g�K3痎���J^��<rͭ�Ư�Q=J�V%��Q0�!�j�|����3��@u�5rVP'�Pl�n�T����~�B���\��N�~��2k� �P]�o����v31��,"o.��D��7�L鐡���������f����N�����B4�,;k����i��xp�V]�<?ݒ����;�@b��Mج�/D�9���C�3P}�[�Li%tLE�2����K��TȜK�o ��������+��@	�"��1?L\�����kf/��I��P步��;���|*�ZV�G�nN���3v�������v������|Tk���T?�>P�c}z�7T��UwU?�)�Si���Zb ��B�������`���q d�F��b����s�,��p:����2|�*pg�a&�^�_BB�wu8���鈒S�n�l=m�m�)6�%����k��)����t5U�/���F�yn�j��ϒ쉠A�k
��fA��Ն�Ɲ��f**�z*Tq�}(Qx}B5{�s"A}M�wY#�#� O��q$Wt���!�s0rV�+���(6�\}��P�{�ۡ� ���f�D���j�,���������=��U��>��K�1R@�>n�9i}����C����jCyY���6a-(Y�A�Ս
μ������K�3�r5�.\$�fƃT�}CP�c���_筜cc�\Jh,B���L���Ɏ�Ґ�$�iN"�1�}�B4��&��NQ%R��/�\��ˍ��I��[�]~��,3��q��o�h(���g�E� �c�Mol��/F� {N��m��f�n�A`8h�W"��WmMPW�`$C>*C���]}�n0��a�wR��H�㨈`0D'��$�_3>n�?�SEkPE�3���<0El�&��b�ɩ���Ɵ���9쁟5?(q6����r��
����v����^o�ח���(gILO�S��Z�k�w|f�pѮ�9�Ś@��Z�XٙT����i,X��$��`�l1�f�����T�m~��w�7���2>@�5x;��M�W�1T�����!	�$�t<��T�Hg�6�Θ!����k�h�rVJ/r���Hr��e�o�/G�bKZ��n������+,g��F@~U.�j!�;$��!Y�}=�յ�TJ;������<�ߜ`�IN�����KH���N}��N��ǥ�-�.3[^w����%b{�s�oU������u#���XJ"��z���^�	�wUbaq�F��O��4���(|�*�vX0z��X�����`ِ����x?	̀�)�����i��$7<�.�D�`������ls�H��.(�*�b����Q��9��gE��N���:�b�_�(+k<#�	3�\��+W��ܧ�n���m&�*J�ұw�>�yb5��Z�Z��	^)��q�7?�E	8���������*�c�  �-砒ߨ��H��8+�4�!�3)�೉3X�(u��.ԋ��y ZN9����Td� 	"]��3���f�%T�7�i��n�IA�t�	�S�^Ј��6�M�ٍh.)�����p��۳Kܞ�P]d�^������t�bK^Z&b�z�o:$/b�`��!.u�'��$���бk	'uI��4S�K(~�o�NZ+�=d�gm������M���t��������n.b\�������D�R����]��́�:�T���3���v8+̄�sfu/�q��x�݅�[ ��W� (u"��'��x�x���G>q�B�c��)/�;
[�'	�<���'���{�UMX���,ϧT��ѱa���-WMvN!2���'�M�ՆMPP�M���Ƽ��v���Ё��}I�*B�GcO��EJ,��)��=F v�3��9���53�+ec<ٹVm��?��ѩ�Ok�sښ� ���'�D)�$U:ji/F|b�r�8Tl���{�"�R�,��XI,�� |���B��WJ�>���4΃��.AC ��iW�t���?�լ�p���y��\�@�s%�%�d
/����ZO�N8_�����[�2� �v���ħ�G� ����y�(�5K�ɫ��7��~��_�۹��iC�?�Cai͐�YbG��Ut����/x/v��Ws�7����f�?������M?c�7�{�l��j%С�Khe�ZBP@�6�5o��$<�1]�Gb���b��A}���V�wM�!��T+�v���9�d�qQX��V�\��!\��/�:� ���ݮ�5�bJ�r蓔��>S�d0�[�^��V���M�U:M0�A?���n��M4"$�Cc'��c�e\��ϝ7�jY~*v�u�ĵ�d��Nt��W� ˽�H�������-r���������0e�L'�	�Δ�)=����j��N�sx`3�r�=6��q,y7���5@�}��3���2������¬���P ';Z�9��j,<���`?]9��NU�i:���w�M�?8������q��03�?N����*���Ͳ���}H;	C<�e

3>�*Q��L�%����?:�&�蠸�p|�3O����wNB,Ln>�O���p��a�E�W7MN�F�GD��8��ʚD��^ҴWK����K��`��W�����	G�:{]x�a��n�+U}I�L����P�vx�+[��:w���@�gp�|��.��%yE�1!Y��;m��B�� �y
('�t(�X��+�ש�x09l�CR:�S�qY8��Ϟ�2�����v�,�L�L�ű��0΁n+v.υ���C��H����aq˂�)����ک�۶���\�ջ�+rxe�+*���jB��L�<�:�x(i�Dr%�.8*���D� ���F8��M	��.*���<Uj���.�6�H��B��\BT��7&1m����DڍO4^�RL!e�I{&�0�"���zu��a0�2�L8?�q?S9U|ϰHf����-CZ���+S(��R�{��{���m�up��-�C,���K~�F��`��Tܘ��	��C�7�f:;g�G�v��Z(�^�� ��	iXnhRE�2��2�q�^󁁰��=��/�ԃw�ׁ\���e����].Es���C(��+E7�D�mP�c��-�����$hó/kc�Q���'�{$M;E��h�{�a�j�:�ş��0��]Y㾼�NB�����r�����\�ƙ���<��������,�CKT���Z��ra��:O�02���hÅyf��^�;���m8Z�.�l��.�Y�����*�cx6\Ы6�R�CJ�6�6����ddJd5W[�J?0�1�X�����A3+>U5mt���Է#�}��Q��e~]�� t��#}JYN4�X�ދ�n%�Y����M{vD��}��S�J�[J��/�b���F~ֆ��x9���<V/Z��ڻC�S��B�=�*��1����=� �3Rzk����
����e�Ԝ�g���䟉CF^��o�ݲ8��{n�v�+H%X�[5~�]�����|
�0�W��K'�A����JU��W�_��w|H��ض�u�MG�u���i~�4�!��9�V��ѐ�aЫ��k�Cf|�x��'�[�4u�ۤU�a����QYO�k��Z���:�p�KW*�|�z7�w�4�a�����-#�>�){Hf�y��&����+fq�_A#�R���Jr[�MJ��B��6o^��AA�����U������s~