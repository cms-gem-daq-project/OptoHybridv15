XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����L�3�Q�t�o����hdL�ֳ���l�ԓ�y�x|��X�;���G��;kҐ(��D��D����t.�Xz��A�����l��B�M.�}%Pk%+;*m���n���,O�d/�=����/Kb�R�X���}�#�� ��"���j����>p���;ѹ�Y�o�W���-'�½^=���a&�`�*� t�SĿVZ�t�Y95<.�KV-t�i�<��y�̫����su 8>ܻ�]�4�@.��
�u�~�V;��v�^���-�(˻AO*A�3�&�Y�'�*�N����DY�O�&w�X���I�r^1��Ǘ �u�%�U��X���$
:b���G�K�ϔ,�;g��9y�GhZˌ���.��
���K��p�[�������&P+b��t�i�M�3,B����m�����\u�](?#�]G�V�.ܟ6�-��9��M�Ej�B���/S��Xs����rr�YA�B��2"��y���Mfܥ��'�k��9Udk3�m�f@�Y��x���!y�A�k�Og�oC<���VӖm�N����L�~n�s��WW��m�v]c�<!�j���a�4�<��#�)uۈH�)JgŨ��T��O��I�*	�Y��ZJ^������4[:�����B�߿��ze(��l�k,����!>4\�p>IL�=R��=��ϩ��P�Y�G
���N�4:�D���M�thŴ�B�h�eRq��O���f#�F	XlxVHYEB    3c8e     900s;n������Q#�V,��z�^�Qx��T��'��R^ <��I�7�8L�P �j1�I�<���/�"���y������� X8�T��?4]��^��n�����jmz�`)VȏRdu�~7���6�q�����AǊ�x�����&=f��ER��������>���H��Ͻ�к��.��L�Qف�~W�W�1�tNC�VX�*p��K5
w�k 9��O�kBo�Ȃg�9���/�PL�&�&�Z�q��}MS~�~�d�b�^�\�����fF��^���j�9�"}07��V9�yO��K0�~#���f2[�����
I{C���R"}�+�� �.vE�A?�ʼ��X@�v���I�_�V�>�M�Nߜڊ�'|� ��R��4�`���xP)�j'�+�;J���?������>�Qh����W�L��R~a�z���tQ��K���������^-�F:�3��}�����gO�l���0�Ռ�!�m���x"����#g�䐾mV�5�Ivm\�7��ye�9��-��@H5�L�E�ض42!�UƌQľt��u>���r���b܈ 07I�VxA#Z�y�d�pYVl��g3Q�������e�'��Y��-4U�a��'�S��z,g���[1��W㙙���L���G���ʟ2T��xjThC%�gvj܁���LK�nI���%9�f�bN��|X���N~�/��o���Q�$/�)�bNcAk�
�|��Do�p�Y��E����%:�[�rv�C��Ҳ���/1�sx�<∰�X\�z\�f �
v/ ���f�M��2#����RbS��0�z��#�u\����M.9���*DR6���?igg҇o������f�	�I��}Zp�5���`c��`,fu��:�e�8_��F=��
z霰> �Bb��-	s�h��� �
ϖW�!�[X��b �,[�\J%�VǪ���b|�蓟��ݯ7"Q+˱��ᶇ|�e9���ʶ���P��)p�i#��a��7,#�Yz��6{ϐx�`UX�@�0�)02ڞi8�c{�D�3`�Qp��{�۳�t*[�م�t������Eο�\��d��QdC)?�_�k�i���Dfxu�E�I�OJ�?�{)Nm9$$�(y�%������I�? �y	'v@�^J>�q��V-�u�Hp�CA���FB�;�>�/��6@C�\n���e�Ԣ�,,�Q���I6i~�к��j����x������W9��S!$�  �-����8�E*��0;��%A���a��!�6��B�3A�)/�Eݸ�\E����T1��?j?�?��� (���=k<�8�щ=��R),��4��E3s��;���M�7[� ���>+G�Z��v*y��V��5�[�T{h�[�:�>3�B�>��q ��62�eګ�t�Ud�K�X�$ G}Ё��}��_b���LR4�q�y#v�$`�}��t�EY��v��{&�Cr|8C�:n��H���'��.�
]�]�D�`������.<����.Ts�0O{ۧ��Ť���-�1	�j�юd�� ��.�l���=�b?��c#ଋ�.L�fV�B/�N�˧4�)H�,+��X�vh�oe=��`�^a��y��o��F�h��	.�oa��k�o^�<�y��f�OO3[Kug����^-��=���k�4��ED*K�C�N�7tu��x�Q3`T��y�xȍ�I���u�Z~�|���Ə�1�4�ړn+mG�����g����-�k�slx�:ȹ��ky�,T� g^�mU�wwRj{
X������m�V�zI���@#u�׊! ۱i=tD�JAdBm���!���n��.R�7�7�ڍ�d_�s�+�\��L��`I�dC� ��v?�����R�ӓ�oL5j�U�]킇�x�{���H]#��^����;���2-\Tj*�I��iTK�i/�ݢ��#���^��9�/V��R"�_`{���,E�h�j�ܷ�{~x�A7�S���INP���z���O�y�D�0��:`+n~��:!װ�G@��D��hYH�����uX�,! �p4\V�U�J7��RV�d�RIC\�����m�OM�a��%������	1���m}-��ɇw��4^�R��l�V�A�{X���cѓ%�&R�n�'zsce�M������#7v���Q��K�c�@7e�l!�X����" �h���Y�5tf?BZ�m�fL�_�����g������:������3+��^`�R)Wt'=�n�