XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3� �8�jb�w,k��DS�a.2�K��HI����SQ�SE7����^hab�J�� �$��j�� 7�8����T�/6�#�h2�%b�O־�W�`o'M���d!6��=�l�R�H���`u��Na

�HM/EUc�@�i oj2�p�rx��&���h���/^��6�S�G\.ݠT?�����	��tb�{[o/]�$y��vTZ�5���m#���M��E{Ү�_"��c��?��_��jEx���I�Ke�>�P��鐽'c�����
�H�a�z��y���o�y<��<E�����Ҝޟ�DV����<��x;��P�55�H�W���.ua�}��v�p<��~"��帎��Lw�m�@�� ��#�ɏ�5�� �����2>E�4I����l��z�Vu�!ZT�&/Xh��2��8�@�ҡ����K&��40��8x��_�����m/�r�%^zw��6Q����OMXFQ=:��Ur��s^�O�����E#��'{�`��[b�/Y�H�����Ix��Yh��
��:�ADMM$�ɖ�P2�f&����`�D�iR��&��E��4c��5�ҾG83�d��̼���wu0j��D�x8{fേR�΅X1����g�n��>>?!(�ao$�z,�qR��R��>>�tB�WlͿ�u3f��i��C�?��YmC]+�`��s9�x�^B�)�g(�b�eܣQ��5৽�vt�������M��Q�_��e��(���ܲXlxVHYEB    312b     7b0�ۦ�%�6�����_�BV#�l�/"�`���'��3�~<��^��(�d�
W״yiK�$ ��{�T�|���r��Ȍ�M�q��/����-�Rw�nO�L�x&ӌ;ǖ�H���
���TO(�s	X)���H�S������?z�Mñ��Z���E^On�"����l���\��ɜN�Y���A��y�k�z�+�@{�;^��cw�M�.��t�QX	p��;:�i�5��+P��u��Į:���Ej�p�B�F(F}]�g��qA��R,jB����*~J������l<�0��'L��+�g;0���q��ev�a���̓�8U �ixx��K}�?s��lHrެf]?z���^"I;E~�����2���;m�{ѩ/ƣ���-Ͻi��7����Z���`%�G;�5%���
�e|:�n"=a�i�����$�0fVɢ���iϕ	�t���)b�7*{xy��EX�S��?K�PH��~�rݡ�r]�˭j�����嫃��"E�O�δ����i06��Pb��.���+z�����)���3�Z�]��� $��֣�K���,��Ю�c����!J�	\�y�.	č�B�)���:���X���8ݓk`�&|l_�y-��&M�����--Fg�M2go��K�$l�I�������JiT�ԏ�5 *|;W�-L�E҈LUI��lT*��ѝ�Mph=�f?a-
]o��pA�rbzo8���s���+��#��d�r*�`oä�3i%�`��v��p�]�\
�	�G�b�:\���}��f��4�v��ֳ�Rr��H�ۭ�nHd�(亽��Yɸ�{�b���)]��G9['H��b��!@Y�_�k��L^�2N��MtY�iھ�.C�o��/�i�]Ȅ���NJ���#�<}��ڴTm+EꎤLt&�b[��_$N*����ٕw5�j�2�t�������d������3�ϙT�%��nÆ]qv��f�Le��� z�Ƽ���Co�й@9y�Z<D�5�o�S��@�.�1l�#�)�_Y�0�y����phQÑ &[!�KT-���Q.
n�FJ].�u�Uc����:�Ӭ��N�ƚk��������]ud�4�,tU3u��F>/�����cjͻJ�H�ؘ.��m�\P5��K�Um���l�f�~�,}ӄ��-��� >�n5����NZ��H�2�e����|t�*ޓ�#,[-�V(͟-����HZ!�!�T�"WlΦ����[�a��Y��~�+�Ѝ�<�ۇ�Y76x~nK����R�S'���th.�v8�|�j��L��� �]�������%l"<�V�\6)��l��6�D�t�O7vCW�<c�&^k���>ۓ��|K�B�(�;�h�����^�2Tw.t�����6����D��v���Z�A�`.��u�)�^�I*�ި���ڃ��K�@�~���/4�y����5�ܖqHp'����U���(��N����֍���㋸)�0$�u�%L����{Niq���T$�ڄM:\�nC��2�>�9�-�A��՚K�>"=uw�T��2Rf�o<,��{��2wB`�g!},x�a���C��m��y�3Mۥ�Hg-���!�mO���s;s����Hy�X��x���s�)����h���0_#����C���f� ���n|Fc�+��E� ;p���&Y4#�!/x�K@�ހ��~Ҁr0ə��kFWK"!?>�׈��\ǳDEE�c�x7��5c��
5��5���>~Ni]���<��P���j�Ќ`�L�&�7iK[����Y���&�߰$��̭[��DK�c�to���j>a��4�3A`�U�{ք�	���4�9fS�ԉ��� ����	�T�sYħ@�R���e���,?����"��h���G+�;	<����B|�Κ.")E~���vw�7JQr��ux���)�GghV4Jc`�Sf�=��tA