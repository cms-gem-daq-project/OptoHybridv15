XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[����z�ݪ�����P�����ǸX,�F��<PR�[�'��'�c;����!
&�8���O����P�P��$�>^R�Q�l�|J���^_��h�������}8���~
v�|�$��Π����?;nP��B�7�a�uz�,f��?���~v���*[��]�h�.a=�1 �|�^�RB"-YT��aF�c�s	'~S��-3�w ��(��"����m�Ӵ0/F��r5�@�aӉ"�T6���L��1h��2[0ܬ}������F�c���r��3�f��|7�u#���V�f]��e�պѸQy]����X~��򩑽�=�
DB����s_�Vx��:F�i������=^/Fh�|'�$���cI�?��"+IIx�+��z4�	�\�x}����&[�1�ߨ�t ���6yoN���{�GF�)ۙj�:E�M�ݒ|��4���,#�(�_7c�@7i�J����i��K��)�Ew�,�u�'%�63�d;��p����7����7C��D�h>�I5�1 �ýU��'G��(~�k7�����e���li����6֬w��Z_L����NO�L�՛�H�JW���-�'�3V���+Nc���$D3lQT��7"u�W�N����pe��a����q���`$��]���y��+"���4���>��B�r�=X���p��賅��E�]�8v9��W��{?Fq7��,������r
0��Ⱦ(��XlxVHYEB     748     310�!&:8e��M�63��3��9plF�g6t��i�C�,�&�幪۠�V�eR�X8�f��9L��ƫ��Ŗ�Y�G�/I�v�c��7[�t'�{o/��b����Z��JsK\}E�G��y�(
!���F�/��:�� �Vx?-[��:�������B �<�𾌱ĤW�R�̊�ݻ��P��g�����#�S��!���{�������zݞRu����馘���G��h���R����QZ���� �k��H�+pS3��Im ��=��5��7��FR."����Ze�l�A:�  �Z7�/$����ȳc{�%Q��Z�R�Ў4�g)q/�46a{C=�AE	 �-�����$�H��U!e�-��{�Vդ�',�z ^�S��F�*�	�Pk���6����Y�7��^060o�r0�Ҧ�3BJ�3�S��b��')�,�?��򤥍��Z�4���U����õ���Ǝc�A�8Ɇ����V��D}܊�{Dbk^�<ə���O�G>@([�d<�ޅW�(��J>�\�PJ�a�+ݚ2�"z3�r`�][����2_ ��������Qg�ςWMoz]����Cf�Y�Wll�zE��F������։8W���J�Q�*�8(����BY�t/���֞�e㑡�#�3�Sde'U�0.�>����6��Ns�θ]ѕ�SY�@;�]�]����@	ҀB�f���W����>2-�s��D=�5�r'�W8�o�y�o�<ݽ��t�)��J�H�F���q���