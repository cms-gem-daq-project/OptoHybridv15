XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�>)���]<!�Jp�T峏���|� M���r�P�vA}2���Ī�#yǴw;��R��>�X<b��w{A�uĨ�=�8#?���Ea���n܅�wfAa���K�m�<H��%[@AUz�]�zL�F��Y�+
3`��o�����h��`!H�2P;��mn�eJ
����K����f�{ĉf �)�=G���bS��A��q�1&�8��D�7�����-�m���u'3 FĿhQfS��-�xsުX���w�bzb�X4����Գ4�g2���ʕ�8��/e�q?�K�	�`>�h$V��=M��S����pL�3f�4qt��������T�o��#{Jڸfm�������٭�	
�ȟ8���к��S�Ǽd�C)���~�{�2L6�"���p�\�H��G�O�|+��^-����(��d�s?J�v���>^�)�%v���3o<��� �/���o�M[d��e�Vˠ�ܨ�R�?�_j1�j�|B�$6���@M%�����H���:���i��Y��$(k[�xC��SLt����г ��pO�]����]��u��}5o�������H&9�bx�.���k;��(f��.��~��j���	���P�=���]�{�!���ί��ArR}E��rK��� vؔ�D�\D� �~U�ꯦ��i��3��/���dO�]����⍁�4{�]I��A�٧���.��bȜV&��T|��
�vlC���1�>J�S�?���kXlxVHYEB    152b     580��-��HZ�-x<�~s��`�Siq�4=����f���0.��D�h. ��i���/��?��D7��
lEf�"G��G_hko����A��\a� ��݇�ڔ�����f���ūsǎ2>���Ӽ���t�L9-���AZ���!*������l��x����
���ۂ��R�Ƿ"�DJ���%	^���U;�� �;_�<S9�y`ݗ��5[�.UC�АyW[c�����9�V��	K�hy̸�T��H�6K�^�jC�Z���[�[w\��i_�>y�W/�fW����4~r�R%�'zB���'�@����Rϟ��lj�6�3�>ٛ��\��??��z,�h���P���,U70:ʭVH�8G�k"�z��fp�Wb�$�����+��/���W@L�N#\hIwB��W`Ap���KTÉ�
�۾�B�����	���߫�*R��i��2�
D\�տj�rII����!�!l[���(F����I�7���8e�^���ʴ��7rZG�#�=���{�g���px���\�Z��b���S�Q���\�(|g$˫��RG�!�+�c6W�5���/��v�C����7	�r�H���.Y�M�����D5��W�dG9��J�UNp�g?�e���8Hg�z���|�4
�w2���
�O V��˦3�DL�M	_��cD>����W˦KV~�_��M!�8�H3�&ϗ%���̚J��v�;�o�3�ew ��G���x&IZ�7�e�$e���)�ͬ��p���ڐ�}g�x�t�}œ*����>m:��Gst{��Xt���-ڇ�3�E"]���j�х~+pK4%e��"�,�AR����8ܝ�*�Ydٷ﹫<~3������f4<4�y&�O�UӞ(Kou?Ӻ�c�����x��8�l~��@(���/��cVI�m�M�o��]-ŞJ�'Fi0�1i*�7^���Jү#� ���޿��#f$^�!������A�~?�O-RhL*{__�� ;i��v/_��/:ѻ4<9��M9�[ϸx�Ñ��~f�4��� ���όU
����vs4��I=���n���3��JDJ���F$7���s�SBCznŬy$�d.u�Q���ݰWx���:�o'��һ&�&�d#�\;�ֈ��}��d�K��LU"��Y�֓pWH��]է�Xa�� 6�ͭn����E������d��(�&�m�n�Yy&��dT����$�6���i:��S���3���MP�:P��8�`�6D�)_ECAbE`�S���̝g�.�{B&�ʜ4���8�8Pj ������i�
�����|E�V���/�����b������y3�	����3��b�G�X\쓙̢+]JJ�hx�?�AL3)V