XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]ЍPNn�fʊ��^�g�W(�+�$�������e	=8�^�<��`��,��4u���lȫ��.43��N}Ƅ[�J���1��Q@������ff��,�p�:�
������A�\���7b��Wƶ*\���DUQ�tT)k��hA�-��u�����?�^�, "w��d��
���͵j�j/K��؟\J]+�LݲXV��`�/��<�5D́��j�|E�W%|u(���xĂ�&��O��H��<��������"��X���Y� �������[!^'>�9��!f"��O
[���+w5}G��i	�u���i�8븥����~ⱷs\�.����x~:��ml������h5��os~�G`�(��i��T���O ��a���9�mN����ό2��uvjƟ�����}�Ns�n�yg奀��:��,k�������K����o/VF�7^	v��߮�M�W{��r�7%�W�k�L����M8x�RRR���l����<]53�n���K(��c�ܱb����Sܠ�h��4��HEk�}7�F�'������@GF�4L��W�%}���@Pw�"tb/.�b'����,j9Dn��˷ͭ� M]KD`�
���s�ϑvj+_Ut�9��-D>������T�E��%)LЩ9�G[_��ڥ�Մ=o�)���aO\��#�.���]@X��M�v�S�oEO�7��cX(*�b�H�D�i�T��7�}�����$��H|�}<1�l�3tQ�Y�*���
���eu�XlxVHYEB    26ec     8e0氰"+k���Jo\6ұ���o��Z�l���z�Yj*�.��n-�Nr#��h*W��+�D�G�4������=�(dYz����a%��٢\�IQ��d�}�w���|dXV�h�?s�����qh��_�c����=�����)Vl]�,M��֟�l����d-��jD�y���M�?X�OtOB��r�8Tl�E�O�F�S>��Ϊ�Gq�+Mظ�c�(�C)\`t���fNF��ݠ�� 	���K�5Ca@ͧ��V�՗����e�<Ѩsc	$��߁��_t>���NX��W/�����$�_�8�G=���>#Q4o�\'���� K���#x��K�Kt�W��$�B�̺���"�酙.��,�zͩ�zR �q�{u�r�����~�&���i���y���O��Ľ��+���4�~��5#��DP�����,3#��G�?}߁����=3dg�B�\�Mm���
C$*�˱` BQ�̚&TϭSڦ�B�Q2iW}�#� ��e5�קT�!;jx;+��8�?� ,hǊ'�.R��D�\N`Rw$2P%+����.b���n��X�e>H� �۵��C�S伵}�h~��|�Sz�JF����n�8�U����y�f;^�f� �[#�=ȗ��f�3��rH���,������h�j������e�˝����]!��oI^·aO�%�(CP5�4h�gW&K?��6__�^��l��#��G�5����hmSeL�;@�;x�;W���J���l� ��l7�@�S�0�] ��#O�[<b�SpO��Y��#\̨�<wᡋ��0eFc�3_�����Kno�˅>������q[`!.}=Z%<8�1����k����J�հ�i�\�M<a���Q��F�i#�,3Һ�o���v�@4�
p\�_^dߋREY�哥���O�Z{&�\�IQ�L��I0Gq_�v�7<��@h~�Y�op�R�I���A����!�]���]+�I������@N�U����)�i��c,A�J�[1.��De��,^���� �[&��;���� 3��H�ֵ�0��w��D�@D'w_l1�ظ�l�<(l��Θ��S���έ-!�i@���µ ��4]B߰��G���9:�׋����^o����]�U�wm09@�t���y���%�q�<a�	}@!�nl�(����7�Z�b_�`��:t�v�{i��E]�}\Б�5�
���aɫ�����L�]�O^�:��+��r9�
.ǫO�Ư����\}W��4}u���S�
c��曋�1�7a��5CК'3
7nI��x��O�D%�kq�ѫ�$^	(@��|։ĳ�����&�۽��['�$P�7�����Lip<�c	�3;�)�u�BQ��ֻ���M6����g�-|���	��m�P��zY��x�c��[�Yua��m~��[[{e�31�{χj@UV��j5�U���������
�oٍebJ�-��j?"\δ�����h��;�O��'��}�s�n��ִ��h��}����W������3̰%�4?��mq����1�sQ��yܧ؇W�}�S����Iz43�]�����c�������iQ�r�#la8�hn��6` �֭���WS9B`/�ַ�E���c�*�i��s��(d=��D�E$�$�$�����4.�,&���S�e=��n�vlI�Ӯe�w͋O0�6[H�s�i��Q}����*x�ߴV0���������=���Ǘ���c�T�8�LC��kօ�~l�L��y>ah`$�u��@I����6����f�&�8v�Td���}nf����~]�	L�e-���)�=��_�G#�1V��* WX�N@�ʙ���T����.I(��sb�!�����B��{0i�d��0^�'Ӎ,ن'�� H	vƙ'^����Bv �����\*�Μ>����?������]�)�%?�FX	q��)wH1�[߿y���,�F�b�"h�p4�ą3��M�
���9�b��{��Ƅۓa>?�R�,���8]�C����#��^��������ٶ��
<��5���h~8%� �'%/�M��H�<�l�Pz�� wt��3�0I[ť���U�����H��Zc�;D�����PP�X�
�q��U��c'���vJ91~�8eIrn�r��\V��������i�ڷ�;h���T����n�H�uO������z;�c��S�ü-*�y~�A=%�\�^��ʏ�i`vĂ����