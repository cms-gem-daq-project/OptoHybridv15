XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������I����Zz���~W3�w>?>�Y��6A�K@�Ő�-�/1���ǄӶBJ�(	��IXW��:�:��{��cm��s�U7�r�,s( ׻ Egh�������X��Ҁ�o�'@��o"�#5������{�Ȑ2jC�K֡��m��2�>�D�X����X�X�ݒ��S3ʵ��\�.6A�m4��=�+�X�1x�(
P����"���+����}A��'>������Yj �р�E<��iQn@�7���;�Bz��F����B���J�?*��/�����[�{���5�:L<�� 8N���E_|N4�%]e\�@C��-/:�_�Eg�W�Y�o9����w��6��$h��7%��j���S�K�o���@���[4�.�`l]�������۔8	h��"��ZK�k���?�� O3%��ݵ4p�W�����VAޢ�@G�@�@f�zٜFj�������_g#��n#���������+#�fR��������f�M�ܶA�\�n�� �U��詪��xrKJ�kD����(Ȍv�>��$db��6����_ᥜ�Z��F8��S:��:1��c�L�- �a9 DU��[�ӋZѝ��*tܱ]����8�<�q����*�I�XGQ�:�O��=�~�w�d�٦�TC�)X�~M#���Ϟͷ����]��9{~C}�/�۴}��ᙄ.�o�ɔ����(��Ϛ�bUES�n���/&�k�OJna����*���ZYqZ�XlxVHYEB    41c2     c40K����0�ӻ��T:��)L�t�����Ɠ �ZE�5U��90<i�=�J���S����ɻ���)��b(b�ew�y���)4
�*���C�9�.V�L�L��"�:��)�)�6d�S�`l���Z�Z53>�D���G�{�B��g���%7�.W�{��*��,K���M�cmw#H���P��5�8/�+5r��7��_D�Z���l�|*�u���$m�i�<�G��ϯ535k `G����4���	�B��O7����B���dŬD|f��	يk�p�� �����ԍG�LY'�hZ��yѼ*�Q�^`T-��֊�D�WŮ�����4��[n�����a"Yj(y�V��D�'�Y[T�nD{9�[\�Z�U�T۬�%L��_eߜd:
pX(���8N�;Q7��ղV����7��fZ�n�(��;gTcm���띋#L})Ij���2�P�l!׻I��ͥ�Y�H7�Ը;r����jrbF�O�K0�S0]�#J���ݾ���׾.���84��Wc��)�����w���3D�/���&L�s��+��nj�e�F�[06�X��ɢe�������m�n0���W��-\qj��y��:m�}�E|��R���kL�$�`�K��fr�Rn�-��ֺ��O�J�;����A�gɗi �E�A}N�t����ƴc�<��O±͖k۬��#����e`���w�к�In��y�>u~����g��bA�Q��>�I-�`�\W�#��*��"*E�Vv��@�=���He��n��� {�R��jv:A�V��h(�<u�=i뮟���wNŢ?����P}1���9q�;�;[Qv��]2���Օ�����W%V�0JҒ�I��W;"�H^�kr�����ZXVۑa6�:�p"3OY�X�
tt�h�#�
BMF��3��y��q?'�lg�?�����z��:�W��Ձ��~ޓo*�ܭ%�l��ӼZb�C�#�8P�@T��d�V�z�V.D��d�:Q<d)Q�"�L�����zlD�����W ��t�$F�"l���=��lȮ�a~�$m������+hu��<`�;dF*͡��1�'8�j(fk�#3Uҷ~0�uEO|�qe]��CC�5�n���>g��+
��h%ry�C��$?�t4C�8��{�-E�ä���"�}/�@��+P�P��Lf���������dLpAN�_k��Ej���M�p<��LZйz�Vףj���A�L�4�Ҡ~sc��lLqpZ�u�4����t�N�=Ѝ���p�Ja�	�S���Lk�Ƌ�]��Ɯ�=]�
����+�~���"7�sI������6UWF�'��>�?��hhn4îQ=]f�*&dX2UFP���V��vc&4M�,��Cս����ǉ�}뻜R�LO	��rP|8�S���Wބa��k�Kb�Ǫ�p�h��s��d��i��A��S�l|	'?}˧#":C	�
�R�X?�/�+��/Q�z�${>���V���W��1o�� �{CG���O�����*�:��sZ�&Ks�s�u����9��2��LȒ23�x��9��НdD�"�l�e�7�kْ�Z�0����s)���`�vE������"f�M��{� %'�o>��8����}M�9�W �k�kJd0#c!��~�!�z,�@^'n��V���}C���M���[䏮�wX(�<R���0ڏi�%�i��{�=��������ox����9������i �@��r�����մ��5;z�Dq�ckwPXE�d�x��4��ʒۜT,���I��dy����il0iR|�a��-����H!j��+gO�d?(f6�?K�1�h��Pa���g+a/?"��J��Ϝ�|�\����l"���x(к�]�N`k��LB�ǹi�	ܢ�39�T0|�y�$f���4�H�'N�
݀�4�MQ��c�A��M��U?
��U"�B#�l���q�Ix8Ȁ{��{��I�o�ÄV��.�n�6������k��ֹG4��T
9�EK���^YBҕ������P��o�x~ �?�[��t�6���IĘE�I�3X�U���pJ������"��B/p�P�O\�^a��E��[��T`�$�0K�:y�C�i�����K���b�aW���a�4����P�8ۉ��(���X<��ǋ�7�	Lj%E8�u=� ݞ 4���pѵ,8�4vw�!��ϑ|�����6l�Sp|I�*] �g�f�[����Z}!�ӋJ+h���~j�ކ �<"�h©t�P:�v'i�x�x��l�ҕ�<L^@��){��1��d�#%��U!^�����I���sBpC]�ӳv=Yr�iE�g3)%ay�L�[m�2M��%e��ڥ�&�$����x��^̈������ݚp�"ҫo�}#��1�W�X68��Wy<���m���&�1���*&fY��*��C�#ĳX�^���#>Ѡo��St��;p�4@��̲�b��WӠ��dJ��&��ؿ��=X�0k���P����89������һ(P�d���1��ї�\��]�m�D#�߾���'!��4�+�ω�:Ci����5����9�Y'�}>5�&���gqg�F1_a�Q����6�O�ĉ��}��_�u�ǎ�	z~�""K��	��,jC���8|87	���	o�А�����k�h�Pֲ�-]p%d��[��%,24l���5>��vSs���ªq���_ J]ln�M�ם� �	�b%�C�D�'�UR����#�#��'F0~�h�v�'��&盙̖�_�*۰]�+�O�7K")�?�;HhƇ��KO`��[�L�
<"X��E2�sN�b�m�ׂ.�-���2I��%�7s9# կ�"�D	��]@�<<� �<?[w��}N��C�����d* N���!v���k�o84���O��A�	J��A_�*��E"{p ?�@yLE�Ų��8���3a���xV�Lg���/f�gub�g�1�ʸ�mj�P�@VP���L�<�vI�{����"�5�p��@�Py��
��D���j3���59pu��nئ�[�3(��� ,0� 8
-s)��