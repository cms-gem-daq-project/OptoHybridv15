XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d=7�r5@����-7��VgW�FG�7����ԥ�~�s��g���,}$�k��:��/�|/o�8ہE���]ɢ#��4S��*��m����ݔ�)R����AhE7�3 ���v���B��8��ZB��wpTr��W�%$7�D�c��kY�
	�UxK���A�sH$u�����ҝ�	/�����N��B5=�T�;\	۰ȶ� p<j��o�;@R-Ǭ<K��6P$I�_T�����hȧ�p���75���z��ԗq+C��u����y}�V�����#��P��gE�3f��q��1�;�w_2cl��V)�S2�L,�%9�(v�p������"@A�`���	J�^��t�ˎw��"	��s���;K1�N��6mj�����4��r���/�'e�R����|L�f�n����=�lb��.&��[!�KF��[	�%nЭu���LNt�~ww�4�DM[^ࡉ����Ў�DG�������p�f���6>
vK�0�m��� �~M��n���\���E`����q��V�T戮��ϙZ���PZ�"��|���mEk��/�"(�m��'�ݲ����W�vC;
Y�EUT����|8�ޥ�>"�U�ɸv�X��1��ҏ�t�G��D�Èp��O��M�ԥ{ϸe/��=��������h�Ĉ�{ⱔ���{+\!a>h��X�S��Wh�H拋�*v��Ê-<C�!72����ll<SS7�T�]G9̺6t*��k�}�Z9ğ7���{D1\2΋<�$=+�XlxVHYEB    5ff4    1040FwfW�I
����A*��R�"H7�L�i�3��a���5j�
���׈auٸ��d/�5c�Hl8p�x)�?0�OOp�X�B�tx��<���Dz���(�J��ڸ:�>pۭ�b@�"7�h�$m@�i&��|j����,U��q�r��v1��������:�͗?=n��н���^r�n������������I	�f����1���<~o�AV���gE�E�ә� õ�-g.��|,�@4,��2"0�jJ��:Q��]�7 �ͬ�c��'�Y����I��̈́+��j'zf��:s�6�(ޅ��iJA-6���9Ƞ#$����o������Pq/�C�M��6��YDp��,�ü�M��~�O����R�b�enD�XN�~�SA�q%��Q����QZ9-�qj���R��5�(���i.�pjMG:\$ѿ�8��/"�Gg҂Е�y�� ���`�;V/�=8q<l�$�O>���@$oM䊬��4]J��E�B�6��Y�����|��4��oJ�t��ߥ���h0�	v!B5L�����[��FM�K�����L=o��j����k�)t1s���Z�o��r;�
�UY�zܐ7�0Bb����,�4}�ǘ���F�9��r�Ѿ��0t#s.��`C��,�U�{< �h��AKƚP����m�{�GW��&���J��a�R�@�)�����k؈����FBȵ�vU�w3��i���gư�#�:毋�)\A��my@���>��G0Y��[��0@ODl?��nc���.������R���F���Xo�������Efg/�bv��.����Ťs��\B�[ϻ�?�F�Q]��b%�n�!����b�K�7�W�{����F���XܶY�I���U`�-��	�l���l]�o`�u�5�P�ڢ�#���-,��7$ۇ��Ͼ�[�����`5[Y���4m��)�k5��,�wmuk�%0�U�o	�tr�CVӾS�
I�,��K!F�V����G*���^��3uX������Y��x��2�߼���{X�����g3V5'q�Ĉ]�s"6J��*�����$���C4(��!��I��ǺD��X|DA�M0�	�Q���<�]^~�ҳ['`f�\y�j�_
�r1�~��?��'�aԶX���"��U2-�x���:? =�Y�F��u��iMAC]��+\t�&�dc����X)�Եo�}���
��Xc��^�I&��6ug���@�ȗ���^q�B��-U*J��g��pj�AV������ށ%�%�h=��3#�e-��}���$�n�m��w�z�m�O��,&�@|�G�l��jZzH�>�$G/�� z��p�g���[�n{�������a#�ak�:����:�҄��+_p�N8SA1^�b���K _>V�7��ޞx������K����{���SI�n�w�D��Ġ{:��i���O��o��C�/1oIN-F�0�9�_9���ί��H孫���X53��� ;�h��qybd��=8g�*�a�s؎5_Sf���v:��T,T�c<�E'�m��{ �~�>(���/ϖ�`o=�j�c��]X��'�F�g�$��y�I�Q���p	{��V{~K�}��*�ę���������iU���m��]>�4�T��p�.֮��N��;��ceF|^�5�T�1o�?lߗ�7pI�ϻi�Y�A�����g&�v�3N��Ԡ�!�MVߐ4��WRB�d��?:롍!�!�|�ueDv�l;]��acQ�������9x=�OMm�|?�3��a��73�\W�KîY�[��[�b(��5>�f,�ieh�'NP�'ڡ�eV���D�R�I,S�K�P�~뮼��|��o�N�bw���=�DO3����S���'I��j@ǝG]��)���/�O	y��ԗ����)���Hj��ւJ��4����������J���ٴ~�����ō$+H84~�g�|^l�v�O�?z��(H���<ŝ�j�eM�����\����N��b���!��P��,���ŏ���X��r-�.r�� M�ok=ɕK���A>/��i_����J�9ˠ�|��^���|���nkgB|���tД�a�f6���Y7�x�<�q��=�ָ�f��H�J�i��S�\�X,C��b+'P4�u&=��}1h�N�6�ݫ���RQ�����m��O3��Ab���
��j��U��PMO�!�`�`|7ۻ�D����~��H�S���M�#��A�k_��#>�\a��u���P?ڰ��k;�uH��L�+�N�@�Yx#�FB�+<������׉��Lc�w%�s�A��]q��5�85���9���-q��vϧ�������\$}�Ư��Vj�LG>����o���1~�;������&O��
��r������7�.v�:x�Ee�e�~��1���I��\Muh���������������K��Md����n|����^3��1��/�ˏ�3�Ni���1B�~���`�]ȣ�h��=|�-��l�3d�k�ՉG�t��0��k��|�1�o�Ĩ!�ˍ�j�t���bZs��� g�DBC?p*R�MxҪ���ew6΃eT���@r�Ի�����Cr�����C/��6�f�'�~��瓐w�ܜ=s]���2�;������� ��%D[O�ʬM����q�j��&_^/����m^�����ӹ��U��������,D�!���=0��84;8Q��y9Fr��j�'��S����Hc8�ϙ�p`� s�k���I�8���8$&�h8{�-��췽k_�x"�X	5�*�.�n��N�B#6����}���ڄǩ�n���q]o3#�wx�wrJ�?[C�_�V=f��eE�
s�V"z��3���_�Ә8�>7�}᧧N�X��u�Zw7�L�W.Ot3G�1��}�9k�WX<��U�8��*7d��W03? Tx^��> <����cu~a����A���R�ܼ(t��ZE��ƈ`èK���:������!����FN�|YF4+R ������[r�2m���'����\t�^<��k����oI�y�Z�5�;p�nUHn�w؈<{����˄�^7�3�#R6=��AT���C��91z�C���^�$����j����WK����"Ư^7�l��puJ�^�5�E����]gU_�C+Z �W� ��m�5�(�⢗ڜ�E���x�pN`F�+%�.��z+��i� #�^i"W��B󽵭G���^��.�?��H�bV+�=�y"�E��[
�����#y��;"��aس b��'єV�֨�Ξg��G�[ܙv� NB����Y�z4�z������.��6 q��6;��b<f�^�����
�r��H	�����_��4'�|.o��O�ł�@R�
�i^�z��]�K>�5�3��ʔ#��.���VMc���Ae���Z1K�b������>I��jL�ԋ�&�u!�Wx�K2�T�]x5��(�ءwh=�.Y���	uC�5N�`4���f���'�S|G7��:T`�]j��W?�")Ei��j��Y8��ȵ��筧�����t�J��`!�[�J��?z�eWn<`^uv!�ș�~�./qtfך��$�N�B��/駋���Y���a�I�&���ӻJE�r�XKe��n�T�E���y;���n�1i0�?	(���7x[Y\"��mP��Jo��G��}r%�����c|�����r��Ԝbe,�H<�D�
�3�qo/u��Ճ��i�u  �֥��)k'x�-��([��$cԬ��
2�4�"��.>&0L~��'Ĉ�t��?�c�|4j�n��Z��\�z��9�ٶ���d{�)��ǒl,$��
BZ���k�R[R9�j��k���)���s��aJ�� �F2��~�w��]�@�r�}��v�����O����Y�Ups�E���+���z���1���X�#-C/�F�����魐)-;&YZ�r��0��&�R�i�����+����[P��8��+���J~ ���g3�)ap�ĩ��w�1t���w�[�;