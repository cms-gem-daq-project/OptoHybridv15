XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.�8տ���iv�i���|CP�w��:�7%F���켭k����;�-S�1���a�g�[�Fô��m��U`�7�z>��jK�4���Q��s�o �QSUJQ_u�K2�A�ˑ�d�;ޣu1���B|�᳔+javNd�^/_�+oxx���$����P M�Į�h3��n� �x��Q�� a���S���1�.�H�0���+~7����_X��/���Hy�S��;�h�!�=�| �w���9k��2���;� ��>\H�Zn�����&�L���=
Rtvz��R/��=))P�%{R�9��ֱb�N@·�k��K��b��K��6�a!4�)�Hܽ �os�x�:�oc��g�x��z2�3*��ܞ�Y������`+e�V��]�����#穌B��<�~�YU���H�~2� �����ߜ4ڇ`���	4#}mÃ�U�Kt4;x�n?J�6�!{-i4Met�@�[����$��~R$"궄x������o`�Ep�s�I��QD�M�t����x�T��բ��D�r�Qϔ~@(a
L���9�{[3�>��'׬t���-oW�d??�P�M}�=0˗E �/��yo)�:apq��NU�{�Q����)g����8���wB���V�٨=�]�֋q�|G�pƦ�<�R���r$E�^��{�Et���?��P2��>P��Hi�;���G��2�^�٦��:���v�kک(�	:�������tI�PW� � h�8����6�s	XlxVHYEB    3246     990{f,f5ǋs�C#�!7����~�H[ç$�ր����r m�Wb'L���,�(3������ݠh 
���G&��%���m�D	b#��d($�����:�����ˋ��x����؛����ˠՍ��ܡ����3�.3k��l�� ���.V�����&Px8�	�r\��v|�r�x��vs�t`�� ���<P�Y2Q'>6�3�N�����f�jc~��2K�9��������#�������Kp`���%s͎(�\��.oe&��[�D�'� ��x��휃�,EK��N$t@z�>�:piذ�Y���A�_�F|�/�к�b.�zZ�o���}ⰳ�>$���14ͤ��Md��٭�O�$�B*��$�����Pj8���9K6��y`6�1?��A�wk~K4Ib a8=�yN.3g�m�>��#[D�a��f����B�g(��)�5�,��Go�ZX��W��a��� �;�:P���n{��B����Ke���B���U�����mq��K��ppe��w��)�aЫT��˙��B� �gb(K��۶䮍�މ��4�/-`w{k�x�k��._~$����R��P�΃��2Z��SW4̕w�ᑭ�$�]H�¬�Q":��SꚂI�F����?�C`�'�q(b}��%a2��PǾ\v�S��j*�3��q J[�s̔��Wڙ9��Y稨n�@�z���B��a�q�,�^/�H٧/�	��a�w�$q�6�Z�>'�N���r	j�����χW�4�2,��$zzuzk��5)����N�'�ۯ�HE��
V/n��=ݳ�I���.����B�˂�gFs��|��>����0k�������zD|���вx�Z	"�=e$J�s@�[O磊)M��څ�}���m��7�P��'�d��{R&E��x����3\�����pzD��W�o�ȹ0�� ��.����LSJ���҆����IJC��K��~�T4�f�wѾ�اz`� ��  �Y4�,�?`�<j�y��
�*#��w�u~'�:�6�!�����VL��-}�G�l�=x.B�r�W\>�=��^�uKgz�m��M/�W������q.:�r£���7�m�30˃� v����D�����h�]�U����t���yl?_�E $�F��<� ���W08�Xtzװ&�mx%F�NQ�3�3�:�'9)Ap����ϲ�%��u���Gצ���>�:a"G^G��	�l�E��ο���0��Ë��Y��>,�+,��IK�����Ϛ�~Qܝ���F~H��i̯��E�:6V�0�wK�JC� C��/lGk:E�D9����V|��t��A��:���Rr����'�G��W�����ݱt�:��I��� �oˠ'����ɽx��l0@�Jeȏ��7{��� KO��7�H(�¼�`�3�R�
��ru:K����7��Bs7� ������2�P&A�	i9KG� �4��0��Aj?���S~�:�z[��|�;�=��[#�_~�fn�'��(��F�dlda�2L�m�~C:��.p�΄H/���Ϩzl��bD��3Y}�ȹM.������4{�r���F��3�g��j��^^vd�8�[d�5�򤔹ڵ�I�i&�>x�ζ�}RI�ܓk4@XjOv�D:���V!M	�sդ�I�ĸC%�P����}v�����q���W�<�K"S�i&0ho8��k/���,�m�m,�����d�Ⱥ�!K��n5���<10�m�՜'�ŋ���P�CO��x(Lɥ��#O2���6�/���`-p��qυ-=F�uy("7߷J�!;G�4�Ak
��υ���z��:jJ䲳nf��|;A�&8��L��mk���)n���ۄ��(�o��}$(��}!&���	<V�vD���2%D��������#�	!�ME%#��\ƫ[U��miW\���p }�t0�fC�F�o�%�/?����j�_��O,UM�J^���DC�~P�~�wU�C��u���I��WL��LM�����=(D��T�p�60{�yC�L�����I�G���Y?CO#'_a��"��V���-�o�:��ڌF᫡ݧ�zz�./��=;�F�Ь�c�L����)dZ��J4��2���`�ڀ V�T��;�� ���#c�1�1͛H�*Hw1@-Gس�K!]sٶp��2?�18��ĕ���L��kތڕ�Y���F�exq��qh�h�ڑ�>'�㺣�<�\���4�5�Eg�N�#��ʔ@a�l�-@d�A�f��1ZN��5�1!�С��͘9�MЁG�6	�q��@:#L8^uu�j�tv���))�PHk�H�C�LC� ��C��p�7C��\���GUdAe�jr�Pz^�f�t"����*Z]p-��Q�