XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Uk�P�00J������������d�7�kF�[��bb�� ��`�Y�����2�,6^��آ=D�
�"�S�`�T���TsESD9�x�����R;���$a�ei�_�`X53U���
^m�fe�c� %+D��
ԝy@̻9�D3��������J�Y�ql|�j�z�6g����@��
�l��O'7�"�~ɠ����pm�U�v�V�M�8 �/a�F-�Z���*�!D�a��z<q�96��ZM$�A&�~�����ًe�c��N������`ٝ�]����;�rf��H7S�":�wx�~�9޵�����|����ሶ�Oޯt23/UGF)ed�p`�̡B����6�~
�4H��ؙ-Z��j-���/v�y
����_�	��k!�hi�=��$��t��/��NwT�i,�]5O�-���bf_���9��RM�����#�dG�Pà��H�� pBDkӛ�6BY(�.w*�F,�8Uy�7�n�T"^�I�mB�2������'���v���D���H8���ŕB�G㢆w��x넙C�hT�0ݐW������;���D��*��S�A���5�2����6>)Z�G�ɂj,�O# ���W�P��`���/��׃���^d=u?"�(Y.j ���o�y��c� ^�7�&)�N�c"[.#�(�2T��ч�x��$��tx���bG�X}��ŉ�Xo�v$G�L�c<�m��T�XlxVHYEB    1620     6e0�ba��\w����s$> Kw����`��E'����eA �`?��d_�x�l�����xs\n��G`��$�������O,��������� �3zg�1��!5]�t���h��|)Qj��N����qR�����e:̿>�����������x֐ 4tm�x�����+��p�p\EZ��>S��*��JiK��!!�Q�/
1�x���K�X����K-�Ȳ�7Kף��9J�ū�Mv��^�%����������~t�;��@�e�t��X,�xH�?F}m�=�b�P[�kO!����u��}&ܽr��(���r�����'��)d(t�S�jv�g�H���x�b>B���M�r�I���H�=�v�y����dJFS������J�ӈ���ؽ.K�oԛ.r��-"�('�nn��Jܡ�*i�|���P�G2�W����x[�f �����B�t9�R�w_�U�&�き��|��l7F:��,�*��0��W�1�]�Hl��nI^�Ғ���!�@�� ���`q����H&�m���F���Z�9� ��@��T�?'#�.KPS3�����Qc��p�_�`1�����e���N��^�]�(1� ����]B����!5-�S}�ӷ��O@�ZF3�Z�~Q��Z";n�y�,��o3�'���.�@ώ��}D��M��*x�l�\�E-z!��V�bV��z0�H\�f�_���Q?!I��/�?�oG{G2E�J�+��ݥ��{7\�5��]�&J;�y��������wrG׏^ȩ���`�E ���[��rk)�BhN ���t�v���s-Y������ǸM��/��h��Ѓ��n�X��,� �E:?�x��'�&���:�d:~5��N���Z��Ql �;K�2-.�������:ж؝�ғXYO�j�`a�k��!߰r9��<���9�!���U��4
�!揺������������K�T���J0)"��.5(�.�]dU���nw{���Wʡ��׹N93�y'pf���x�ȃcGP�M��Ӗ}���8���T쓰�*���U�u1v���i&�O�W��˄M�NI��J��<sG����Y�0�������fl���gD�р���*�rv''؛�ˍ���bP�$F^��r�T�hxY�!{��1�wz�����B(�{OQ`��#{��6���Ze7o���?�uf�P��+Y�Y�C:��e���sf(�l��:r(��-��.�V�~O�ˋ������ےG�o���Y!wEh�wh*ʸp�0����wB[��$S��=?��[;p6�0�Қnq���������M��NG�J��C�.�ʑ���W[�t�nrF"#��1�墨F�39�ӌ����M�.�nǆ������m>=�^�;���5v���Z�<���A��8"9�h��M�=V�q��h9ƁmQ��f /	����:W�P�)yegiӝ8Ub<sJլ{^��̠�~ˊ�Az�욋��*���.�=�2�?��"���Dic�*�w�-�2|g�o#d�$�52�c���E�n��+8����N���mÍ��Fl�S���ِ�S��8�E�>p���~:�[�2,q�s!�� ����U�`�L�.a	�y2�(�t�ڌn|r%e9����;L�o�+=��ShHm�bJJ�^�0�}��6l���v����qdqw��>æ\�4?X|���[��~�$�s֊M��:�S�o