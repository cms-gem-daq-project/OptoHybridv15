XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��tG�PE�Co����2Oq�G��enBQ�Wtc���)���C�{Zҥf��_se��-��@W��ЧS��5���R�T��].p��x.j�����PW&�ӧ&���P��%��`���wz��ݮ��R���������_����d���Ry�ƿ�=�	I��OYX����=Y��Ak��CL�LĬ��/vV�A���lſu�]����=S?:(G?	�}kY�6Jњ"ė�j���7���1�EB�G����ڍ�Ɇ�/�ɂМ��"+���ʅ���%˺Wb봤D/��\��v���nzsv�ҁ� e��j(.�<�,�%�|>��	��2.��횡m�a���q�K�(�4�``;k)��!%~��c�H���l߅\OB�Ǳa1��ϯ �l$1���&0��a��
r��1
��o�f�-��q���P���0��G/d�Ǭ桲~w�9�6
�6/\�EiN@/:��IcZ�)���guׯ���Ϳ���!AYhK>D����R�-u2=e�:��0�ˠ'ʕv��8+�?�U��J+A�ߑWl+i7[J���iڷF���h��qv���q�+� ��I��+R�qi�Q��R`��Оe�	=l��z}��1±Spo���<�t��M$�����x
�\F������ě��"��I�u�kd0HO��@���p��뛢�qZJU_�u�-��{{�{�8=��K"M�OJ���g��l&]&ڡϙq���ϩ<�	S��L�M�UWf�XlxVHYEB    41be     c40K����]�A�zh��7/�8�A���
Lq�x�|�R���qA��S~�J�,�T�h�B
�鯁w2��-r�}>Rz`��ꎊ��bؠ����%����o*��R'.õ{�� ��z��~jaD��櫰��0�����̱��E���N'r�VY2��}���m�U��Ց`�Z����H���8�$� HEj� �����2��*l��e �*��[M���k��A!�ED���.@c~�ۋ�6��,'�N#��G���~%�C���П�wh���.����VB7L�V��JPy���E$�ڞ�o�J�D���3]2���>0FP=b��к畒no�3w�i�ƿ��	)�!t�l[�3��8����0����>�&4���|�$0�^�&�OF��z��r0�G��[`PG�}���*b&Iq��B_���?򢾟\��|H�{m�*k���M0��S�<;k�wO�&S_���pZ�Ɖr�u1I@ ��a���-J��H����7��?��s^��޴	)dL2���+���ޚ��*�[ <����[�]�b�����\܈����M2n��}�:���d_�5�D�B$@�}5�ɐ�0ͣUG@C�<�0�ѓ>Z��܂�8��Ŵ' �e����趗���2�9��V~��}�y#Et
s����8%s�R*�\Z�l�N�,	�U���F�&�Q��C�\ �z�d����}.F���A���R�ֆ�9<.�/�NX}1�Ƽ�ݶ�����A����ߖ�nz�R�����xǣ(��ѩ��4Bֵ��0�1,�|�����)���c��%�
`Y�M���y";�KG�Ƈ��o�ܥ���dELL�]�B���|�9I�Ь��'Z:��{ *�dӐ�
Q��x[_�#���%���-ᴣ�6�!��%���4Dζ��P1�:�x��6¹O8�ڂ�����V�4b�
=�Up#^R	wdab~�_sB͢#G�J���C;���?`u&�ge�ŏBu� ���}�3�؉��?�u'{ɡ躞)��3�N/�v1�:�/zms�W�uSXЁki53���D�@eP/�`~��+40*�X((�d�Z���-:������א�yH[0�pc��7�o���zbBji4���(@��.�<��]�I��\�~D)$��`�X�e;��i&=;$�lg�㭛��n���'�y��Sسb�����2;4&�C5O^�08�糵�����v��׷m0LT%�e+^ ����w�;�[נPያ��WY�T�����K'7���l]����#��[�dp�#��.������v�)������zۤ��rks�{;��l푳�]��y��%L���C+5�^L
�>4��U��p�W��/��9���ރD�j��]��P���b����*�fX*��jC�o�ZAE����m?5}�I����l>�Zw��%"?��iMjA�n0��@i#��"�>�DA�������2c3�?c�����ٳ����CԪW��j4I��PCA5 ��XFQH�FF5=\�q�ܷfz����\�=�o,����p����''���E�8n�����{N��Ӈ��&���^*}���^'ܠ�7��S��~sX�b�F�D�:�h{�|ڑ�m�>|�#B���ĳy�
 )s��PJ��]FŮ��6YB� 	G >xoE��nS�@�\pc%a�����2�˛ݻ�2�"7��c�Ł)_pCN��iO��:N<>��j�R����D����dw�6�_:'��}�е~�z��l���<��{ۙ��Sż������\����T	%�0l��e�֙�*0���\
�Y�i]��ΫS#?�<�B���,*�	I�Y+����v�-��;ZH|g	?n-�X���n��y���GZ��XB@�`m�&��Vr
�x���Şx*�bٜ�����v�%U�o`�N̶-`�J�E��.� �A�b��-ևX���µ��vn,��EE�OC���b����l���P#va�HoׄP�8�a��Q�ٰ|���� ��ȸǵR.�,U�����Y��f���L%%")�>��r�b�!��|#f�#�z_�%b�@�Z�3�H��r�c�D�C���������'X��X�]���߹1IGG�'��-�6�G8@	�ؑF,�JԷI��5= I���I}��5%��u:�ݭ�����1�@o OPZ3�N3���|��ZU�K%��*{Θ�:Ͼ\t5��@ϋ>P(�|�~dyǡ3jSl�f<���p�#P�Q|-|��a��,$�lӃ��V�>�ya%�ೂU�;�f���)�뽼�N�o�;��~����=M���f=�����,�a�����������.�3z�Z�U��Y	�f�*�܌e+m��r+'U��ە]�kg���0����=��af��t��N�e��Z����VY.5Ϳ����Dɱ�M� ����~+���B�J�c+��I��CN�3F�ݜ
�TD����`��� P�-�1��3+�P��@�X�I
�<���ć�Y��k9"��{�@��J8ԕZ�~��vǨ�CG0N���@�ģ�aU��l�"Dq��j��C�^\>�8�co�J�`�|Ӣ(���q����sG.�y��3��'�_ W���-*��s�,d�^�e!���H�|a�c¶߄�X&j�_ �^�K�A��{���n�kP����Jţ΅#�ؔJ�u~��{�OѮJ�ŭ�H�	�.p�ۥ�2�u8�r�ېD�S���->E�<%!L��"�e?�V�':X2�GӁ)Rd�;��k���Q�yPk.��lG���8�C+���&^1��~é�6ܶ�Ky�(Y�I�s�*�I��H"B��'�%M���Pn��&�f�!���f��8��R{�A9�.��Z �#F'@�b�^ߢ�
��bV�CK^�}�=a�g�'|�i*��úsz�Ѣ��?�}�< ����[X���"�_�i�Ƅ�TG�*���.�س�A.��^h�A�.��ʆu{��\��B�r�A`�
!�����-Ͽ� � ��$�^���{pb���8�-�J^�Ҕ�%�P\��3%\��B