XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����[�D-��=�^�6��Ֆ`�B�G�$d�-?奭�s��(����us(�ުC������9TT�|s~�8CB �{�ld�W� 
^O�Cw!'�����\�.���n���-2���y�18<���ٮ�F��T�He�hYCa��#Z�l�|�r�L=H^�ӕ�2�HެBƶ�<\�*���m��L}a_�WҘ�r�����O��-�]B���߽�ţ�E@��t'nŔ��G��OsMu�g�����x$�ݿ���J;�T~������'җ�ۈ���h�G� V
�����Un�'!e��Ƥ���0j_D�eFpd����Ә;�HC���������&ܕ��t�695�F��M� /B6/@E����䳌�M}�6Et8�_=�pt��E��\�h��	�5�	�5z���q��ZV>0���ZJ�ݑ	���D�'���F��K��mE�	ϗ�&˽IL�,���l��	d�
4Cv��e�1&T"-c%6^G;)������?��}�׎���B���l:�ҬdA�^��Du��T��C��4 ��]��>rTr%�_J����&�?�כj�:R��%��̽�������b�F�ƹ�x6�i(�;l�	��I�=��(�6H�j �Y�!@��7��
�Y|�<�uB�6L֙=6�t�J��6�gJ�}^vHNȪ��E�bƉq�G��'�XUCɧ�:p�N���hS<2�*��d�&��A����N��p�������t �|���u��mXlxVHYEB    152e     580�X�CaODVٿ��K�����%<7
��Dv>���@��Tܚ���J�y���F����O���Nw�����6��>L~hs�W�=K����l������<���Mdޭ��6q��9�H��{Un�!U�[V\�j������l�%m�x<z�|�?w���ۅH Ҧ�i�	϶?�T�0C�X�=R����%��"OI��ٰ�%��ϰ�n/�Tz6ڎOs�%
?��R7uL��|��.�U��ҿ�����\��݊g��$��<Tއ�d�j��t=M�$�Ej����g�̓���TU�w�p�Icu�Y ���D�N��%%�vL���"A��v�"b5�6tTՀ��ek�ʳ#�$pD��t�S�M����(#y"�]�3)q�?G�4.�̄�s6�,t�_�� W	$��{��Hj�_���"��H^^���d *1�.��P;������G�G�nV�Zk�=�4��~� n�4�#�u�]*�?:Ccsl�g�gt���O�Xұ;�wn�`I�����o&�<�-���Pmp'���5����v>`0όV@4Ϥs!	|�$��,�q�� ���K5S2��8��LA�3�v���1�|��ރG��c��$�~�i$h�qW&v�`ɲg�_�cOh��I�x<�/�2qZY-�I���c��*�-��}l���s��V��N��{Y�w��k2�2[YCN"{7j�@Qc'"�e�CWٽ,�ե�%�����Ep��PWt��ͽ���a�Tfd��p�~��i��4
�G��l�q���E������}*�z�:�d j��a����h/�8��9W\)#�5��U!��	��a�	0g����G(ii�4	Ǉ��<M�}0���],�c��0dKT��<�uN4���{��[��ڜmc��qQ9�$��N,!��<��cVl�4��Qq/{�$wT-r��R�|�HT�y������"	D谒����t�.��s��-h��c���3ƽ}��0�v���z�Zҕ�~u�
y-֏rه˵?�d�¬��s�qr5ۇ?n��\x�$t[t:�ZNe�c�P'��{"�a��`<[\��0>�h�h�����t�Vy���72���I��o%�ZoU���=��F� �4t�>�TY$�m_�W2Ti'X���e�~�zķ������m�d�.@'��7=���x,��������#Ee�M�s�"�̝�*�?_ʱ=_�a�&5����v��(b�yMn��P��(TT�ĢX �+:ҷ��f󂥻e��~	w=���M�p���pʕ��K0�c ��g_ӛ���W���dB��2�n����5�Y�=��&�H���jv���U*g��>�s��^j?����2��Ԍ9�l9����/:��iey��9/RrUMeL� �