XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��YK_^V�B�~�pfkSH�0��~�+��c\�����s�^ˋ��:��MU3͟�}��>���aylӃw`T��������ƄoZ�2b�ۮw�Ο�2d�*U�ޯ���q|��Tm[*R�����%pk��w�^�Fx7�J%��#,p�d��,��,.��[S&-FPU�	� 25g-D��i��`�#Zx�ޜ	�U-����^׈�&��ӘR-)� �ez�&�,w[�9,m������ٮ��~4y�E���6���xyOV:aaO$0���\��� ��w� ��=�c��G}�`kQ�K���ߠ"Pl�$7[sz]�� ��Z�Gn#6]#-�_��+�gי�PcHV�۞�����ڹxl��ɜ�,���x��u�-����¨��� ��;痽�z��c�����"��x{]�1Z����al9<5u+�����$R���br�u-0��m���X�r���TêyPQVC[Op�=�ê�M��0�&��p��<�+���?�@>!���S�D|2�\�t�|9�Kǒ�R;]*��B�]��u��0%�4 G�H	}�S�� ] ��; kUK�V���=m)�̪!��� �u��;�!�J��3�������uIP�;��9����>d��" g���nd�����J�ވ�$�i#ړ�A��P/Sw?i�� ��Q�a�Ҝ�9���(�#m���Fzo�fn'�;�ԴA���+��c|Y߹�:!^�hK�d� �W<�Y�m���U�����"\6��XlxVHYEB    11ef     540f�fn"�dY�2������U���1=�@�B��m�2 ���<��[�y���G�cY2�� p-F�����ˬ���8���0�Ē+���>�����7����n�/�X��mBu��֍�>rtKJ�S�e����=,*��݊��+p����Z�zNVn�kjʃ�Bo����}�N�\kM��=�}�\��ݩ�����`�%5#4�c5�Y�o�A��8(���b�i�#W���"��vf����2�Q�7C0����R P��S(aa��x�"P#�mc��Ԫ�����<�4G^�{B�]����N-"��|�׏�����>�������&6�M�"����zk�먯��vL� �Q��i}i�]�/(�l��gv�sVmYs��L��`%��R��7Ŕ�Y�!� ���pt�=%@�CIw2`�~��*
P|�ו�5Vo��O@$���4,d�+}�_*1�ާ�U����[ѕ��K㓨��E����l +;f�:� �ԍG���g=u��:��R?~�{d)޶`/��ҥrsf	<�?�xl���ݸ�~L����U� �h�Y�e�!9>wӾ= uP�߂�9�bz�>Ͱ�Bx�Q
�W8��|G�A�������I*�%g� ��7�R���6�w�乣C��4Yr��QAu��5��:��1��W𿫚p�"y���ˉu���F��Dtv���Sڟ��i�����m���a���aEA/0��8��;��O��}�n�}��(��<5��Wp<������<$���V�ז&�|1�>d=�a�"��LP��"�B��Ԁ�raN��<�9L�G�������e����YDŜ��*I�0{��	-e�Nq0P3��~=FE����sj����=ۡw�b�(�LNL��;�Bv��킇�+�����Z�>��O�[ت�NW��﬍�I�@	� ��za�Ш�.m1p?�\��5���Ԫ4ߥ��S?Wd��K�
�p��c��]q�MgN(�[T�=W���oe �s'���iWqi�G�,MP����k���� �ej��B�2�#&�J+�GӒ�ϑ��i��bm��FՃ�^�ڛfG�ok�^�j�-:v�wA�����PoF�6���-��wpS���G#�(kU��z۴_
���3�+�~���Ɣ�������1���h��:1�y��0�����oxa�i'�И��hhm���+,�G(X�K�jނ��� ��VDic���r�5!�L�b���I� ��6e�'�)�3u�V5?1+7rpS}b�?9�"H6�q\�e&F/b�ÛE-Ϧ�U/7ߌ
�$��A�b9��*� qB��GjIR����cK�