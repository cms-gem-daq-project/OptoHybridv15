XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oXȗu%A�|u���q�)I/y\��*��_�����z�B��t������"w�=N h:1�ȿ٦��1
�X@�,ؗ���/Ûa�C�
&�E�F��@��5B���+��Y���*��:H0ZS-YS�6���a[�zbGε��G	�\�Y곫�SX	�F$���+�2=W���L������%&��)�aε����&!��$);�^5�&f��2�H��n�g��c��m�g:�+a��|:�%a>�������Y��GH]�����Rl�ծ��UFb3��(4ӷ?p�R�B�/�)������}���߯�!���Z���t1�]+�Q:	>��S9^A�G�g�gmi���9¶mRە�G�CwRW|ǀ���j١e�	!II]/�WX�_�y;Kt��l��a�D͢�0�X^���I����%��F\��z�+"Q]a�V��u��sY��VˤwfQ���'�ڶ��$
�.�]�
�6%�&�R�a X�2ز�Qy$8��{H�.��d#�w���L�)��%��i9d�#g|r��^�E�e��y�l�d��]qZ��d�o�[p���G�3  ��h�c�B�G�B}�kz��(?��Np�J�ￊ:_��.k^�����Ց���2���e�fg���0R��Ҽ�;ٌ$�Bldӈf:�cL�L��d-��ny���]��iJ�7c�����U�T%4G���HAt:"�^υ��%~v
���m�1(�Yr�����ަ����XlxVHYEB    a354    18907�O)^��c��,E⫠�4����M��
����o:�����;4xj,����Oǹ	�f�i��z��Y}�)uOZ��"3�҂����rw�[8YU���8��+A�(��sVI��{�a�4�cN!��ɻ�'ɸ��9���A���̄��!��e�qL���AU��e�Y�Db3�ߍ,0IJ�ơ��H��R���Q"�c��א�,��R�����G��l�ˬ�*^�3Y�6q�v�/"gw�=f�NH�m�~(<��X�k�V/F�2p?s��=���5WYN��� �2����>*QQ�����lK�]��j�EА��kgO�!��q�H���-SR�+zq����ě�GЧvҁ��ᢢ�Sx#I��/���!��y@�(��I�ɮjH)!�l��ܑ%_p��P__ۡ�� ���h/]{��"ǶƦ/Mk\�ӯR+�~@�����������0r&%D$��˼��_W�{q�:F�Kx:|)��a;�{d{�[�=�$�RkEA��j}�G7m�e;�(0��U�+
�#�p��Y<:�����Q�1�� ���U�u�{]�߉����'C�:o��\@U0���z�C/x��ՀV�D%�ɺw�<~+ �i(C6��]�:���!��}\���|I�����^*&gL�n��w���������%�e��Ŝ�v�
���5ݡ�q��� V�ɞ +�ƴl��"ίe|���0��g�N����>����Z���p/��o�fm�6�7���zi�#lPI����`+��5*�����yӎ�{׾���o���m�(����9�F�A�j�m.ɐ�=����m���~Q-����䐕�H�a~����]����U�I	�����b�W}� 1;�+�(0���(��sԖ�����D��v'�=K��y������pr������/~����=��S �8b���N.�b7�[x���VS�8&�f�5���1���	��CE�}# ���FD��1h�:����N*~.���l�� ���5`�ۯp�l��4���QFG'br�9��9<��K$跤�s㜗�ca��3~����_�j~��RJ\y��O���S^����t��
��t���Т�>U�"��^�]�� �i>F���?��,�s��E�!ж<�qڻ��6	��3�Q.�T�ȳ��+�D��e���f䣟�E%!�0>.N�:��Js���=d�UP�:!�֮?�%n��3(�2�����W3=^4��PǿKN��e��&�`�ڐ��z�z$���,]G�q}�H݃��zC���	kS�ON�S+	5�Q�G^�"3ejΥ;� ���r���P#5�*E[27�7
V�I��jÛ��U�k��Ѥh�P�"	*��3��ct�Vݤ�n:K]�����v� [���پ�8��a�em<^�O|K��=8��D \�fw��u�&9 *N�����_>ݔ3�{�9�]����O���.��#��{�W��=+�1�c�Q��o���]3�l��k��7����Ռ�;��,���ڡ��V��8��|���cTb�9�P��cF�z��~�J��HT���;�k�2jh�>��w1�;�c(�l�*�1�T�"Ie:�I�O���#�ez��q��pX��;�u���^�є��p�4�d��g�Y�C�u9�[1	���է��)߰k8�*��Fj͛ �}Cc�)�܅py��Q)�������*`�λ#�o�?i��o�H����Y�<��&��Hn;�8?�H����6��\D~��lP��P��d�����$ � �`a�y&�� ������#V5��.�i�����`��X�D$b��i� p�S��u
��E�UW+��"4��D�@���)!�d`�����|g eff05�,�!��h��0�ry�5I;s�Bf�)�P���x���
�rM9�^��5��/z+m3,�Ԑ��p���W�����
�{�4O���A|.�C��m�pg����V�k)<0���bP3�)G�ζ�g�~�?��XP���u.>W�K�o�-�e���a&I��,9��>�r_����WF#�x�q�7���VL�r%>��%>�A����D@*��0�\#`�l`F����B"�R��Z�'�u��5�K�.�|��NHR��K�-��b���CN���ց�`<�W�e�S]v�Ȅmd��|&�}��)��!�`�M��ԝ���v�=8+�!4#+�k��(�JG�Kf�ܥ.AU��,�rK��ί�)�3U�Q3\��NOd����)�j�aY�5o����T�	֜�1��$]�k6�,��k�?z���>T�r�*��@$�W���~[�$V�B�Bͳ��NCtǁJ?)�C�u�O�JF���.����>َ�e	���eTx�^��Y �c��#5���nS�M����,�̓�]X�e�P�B$�GP�Ҁ� L�?`M����.	��!��L��;�l�����hZ�*}�$�����jn��&b���^��q�^���dey?�E՘�q��ԕ���$l��ּ��ґ1㲗@%�eXl���7p�o�d��&��Z�k*��Vҡ}�(/��;v4�Kt�j}��`��^T�B�����E�$]w�Q���$�\���'D��a����A}����v�ݭ��s%�v�R�]r���7K��-�TYo�h�g��2�!�|���ǀ&هe��Y���PJ4y#�ybkQ˫j��0>om�����4�0=�H]yC@�]@�=��r�%����n���ڐ�NP@h��jș�TN���D1���t�ǅu4�z8*A�T��H�1����>=��XK4�hV��[B �܀hn�r���ttyϖ����7��W�C��['5�O ��D�wsE�_���W�����/� l��Aa��K�"��:��ïh	v��l�z������jR�;�]������0?�}�/ ���t-"�!�t�1�8�IVFX����&�ZW*x��UiX��N>ɒ�f��1;����#�b������6��� ȝQ�	�ĝU��`'<b�|	��Ӗ�� ���Ոz�P��_�N��j}6���_�����%�6K�I�.���M=�Ŀ8ݦ�[��1��%�lς;�^��A�X����e>`��+l�}q���w�rcZ��<oڡ�%���h��������D���	��a��Oו��Ly�����ws	N �Ԧ:2i�؍�!����� ߨ�-o~"~�1����T��|m�Pi����d��2��Qe"���A�aN5�%����`�H?*�Ƨ &R ���h�K���_������uI�ܪ��� #8�.)�!�f��D`�f�Jm����e�4���4��s�;�PH���4�/K�F���בh��F�W�;�%
9����A�N��Ϝn��C����}�a�x�~zz�KBA𡚡��S�<:K�p�=�9V�Bx7"^u(�$�����&_u�R���ϢF��J�Otz����&�]:1J�����N�51�/R?zIW�u���C]�+�վ��%4a�Z��ϔf Z�Ӕ�Q��@�j!\���4D�y��Z�6ii��aq6k@5�cy�S���K�	wT$�i@o;�*��:��p��JPf��90����4�3�7�BP��`�o2����q{RQ�\p�b���u�k�?E��I@��{~�m&�Mq��v_�[ҧ`�C��=.�C5ŌT©�X��5`;L��x��=������-�=u��B\�΂�G<0�y��,�����YS�O=J���/�������[�=!P�1X �Ʒb�k<'����r�<`m� 0����oNI�:$�9�qV�ɰx\��I���DY�86%�'Q���M���|��Y�ʠ� �6��*H�ɠ �%$�_�SV�B
�IӞi��H�|֟���?��CM�u�ǖ��^�m��B{�O�x;?�ʪŨ����	K������;�D��J���8n ��b�E��I�-����aa���)18�$���j3N���J~fa��m��ļ�;����	0����ւ��nG�|#��6,FQm�o�tw��Wo�(z���Z��|̦u�
gqP��ܢ6�3���]"��pջ!{�듲��YE��H�Y��#��(`�Ъ^L35��b��� ЊhVB�EF*d^|��?��7��
D`F������z�����({�Tڅ1,��K"��4�PN��rL��/�}��+lc(#yt�0 \y*�'�o2���GP���ő&��u��e�,�W�}
�ƇI���t��¨�ߕ=���p] ��5���(=��zv��Cs6���%0iqe@�R��QM �����$�70��[c��$r�U�F��#u����D �*���T��c��Q��Y���ڛ���Z�_�J�w"�*��gY/H%P�e�)�MՊ��BN)�sr%��!��� ��{��6�ps�_:ky��傪,.	t�c������q{�Ņ�����0z��!��W&b,& ���pA��X\�^���(x���c/#N�T �q*��˘�B�69�I�H�b�x	��kw!��WCP��"?�����V�T�b;�v�ʲҸ���L�Y��P�Y$e�\ �/8$G ��P��d��Ҙ�NN{�~���>v��J����a��x�k�t�|�!]Z�Y��!܍:(j���ƖU�n��0j��/b�����r�l�����Kv�>=����j�������L޹�S�}h4K`������z:��6�,�Ի� ���|LMr�ҩ�}�<iz���n���;��:&�:�*��u*n�|4�0����Q�b�)���>���Ӽ��|��u�2-�e�[M\�/]��*�}+1��>�1W��	Qf痟��U��b(���6����.�8]��i]f�"����?c���&�&��&���T��-������~Lw��S:��bC��	 ,D����]%G�Pp:O���|9��O�	�Q��>l p�$˛c�)��[@ݼG��-�g�(���L�� ���ώ;�y��:�9G4���К ���G{���5��zwT��llӟ��^�c=��<�|��֕�?_��T�����S	����H�>kD���% �C��^�<��#��3�{/��/��Tiv����� ��b\�-�Re3�]�Q��\=�STV�O�r�i�֍[���d��~�z���rcS���ك������2Rr-#���q��Y��U��w5�=�y�ˆ�ܨw~�s����yF��W���^L�d������}�fƻ
��@G>���â��WfW� |�RW@������ ���e���%�9���s��"�VA�����K�͆�M����C��tB��� �vp�~}�$�Ws����E�x��8>ƒ��f�<�ZR�d�m�AA����F����<�d��2
2�*�_��֧7�*��}�DnQ�����4��oH<q�[n	����о�(�+�6>#��퍳�S�P��
fʮɩȤ5A�P���u	��r�X���1v�BsK�K������3�'!��8�%�h�@n���l|Jz�[�)M���7�˴���Й��K�7P�9��!xG�׀��v�؆�ߌIw�4G�9�����mMz�y�-�_|TChЃkb!�|i�믞pn�'�9C��R�qso�$� 5�<n���]��΅k�DR<^����h;ZfRzoh��c,%���4S�4�恞�["E���fOe�I�a���*&�%	lB�XTH*ԇ�6�_d~y�J�KU����P�U��jY��U�q���+9;@�<��i}]0�Ҍ�,�L튾=�$�W��Mt,z���v?��5;���R���wp�֜��|�3y�#�ɂ �1�c�V���;u���o ���^JU�w�+���܈"�4�a �\c�%U�,�ڭ&h�M�k����o�h�+5���4�>
��钦N����JeA���!}d�w�`8��p�=�:�_�': �p�I� w���X��%���a�*N�A,�$�0T:\��JT��t�ao5z�r'���>�u{�n�B��{����K���ڐn�zh�N.L�d\� �˅�'�~q��}�,z�;f?/��k�1X3Bq�T���ɱ˦���F��.6�{�t@�(�xiT��
dhl@5p�㥇����P��ڔu�{+/�OE�=__wC@Z�