XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=Mrn��n�3��/~�v�,�\�l��Ǯ!xZ%?��E۠~���sԩ�܆J무�P�1������Q3?Ɍ?�Ksi"%o�|߳�E,�Vi��\���Li�6;�t����滗��w��E��<VV�t��l|�l�8�s�[m�a��R���9a��(��m�b��h���nR �ݿ��ςǢ��*�����s�Q������"W�^��[��*^CȜ�DMm��_�����3������{��9VDب�#�፲���L4.�\� �N�c��|T�<̧6��w��Uj�l!īq'��Yg��H��5��,b��: ��(f(!�?�����;>7$A�y����G/Ms��q�'�3rJT�:�:i�S��曩�L�Ƨ �Ӑ�#>�%بkW���L;ϩ���i_l=U��'�u���F�t)��Z����d��O� �9d�2�b����Ӣ�3߅������fzdJ�_�S.!THcyڟu,�3�4�V���lR	��B�� �f�.�D��#�2�F{��nI�s�X�0��0�X�HM��;2Ym�^����NV(QR�;����jk�>��ܶ������X��n�D�X~F#��	9���M�	�����d¢���5�mXc!M�ց�k�B���'������<�_��'*�8���4�Pd,�m�����Q�e��,͢���N5������Xp
�|�7
&�"�=��s�v�#���!x3:�`S$AqXlxVHYEB    1578     5a0h��x_��zÏ4WA @�l���W.{�Dr��VEa�C�Y���zh����v>����iM�G�'^�[1���r�x�5k �%�Yj�* ��<h����x��(f��������P�� +�@�̌*j�����Lb�ut}Ra8F�H(���^ R�lrފ5�������~/����O�� ���u4�aw��"����L�����^�Rk1�KwB�7H�^"�Q�M]�Um�L}D��6�%��f0��L���"5y#F�]�{�T)(O{�v�9��������m�25z$)�<����(R%xO��a�\��8ۊa��3��Z���-�<�@"�1�����wj��NBK&yS�D���e�|U��5�^�\Q��;� ���m�ψ�gǘ~t'!$]f��*A���nM���v�*;���h��]�]��vV��:r��>B��xy�D���7O4�ʓ,6�ϵ�M�l}JZ3�q&b��G\�uN�H7)�|T-�K�#`�Y5m'I�"�UK��ːl��kNk�k���z`xL��9�_�PF��㯂�lx�^�4@�%(�����B]`��XV�#U�r�˘��Ds&��k���#��^�.��#��M����u�>���7�uK�0s�lII~�Ӈ#�[!1�,��c6|���PSl-s����r�l�R���N?8���·\ �4����I��mΨ���_��,iEn1b���j��B���9�^Ʉ���(�֍W�aa�C��[L6Q���荄��ݽɭJ�+�fO@c��δ8�*T|���Gͭ h�
d�� �a�0K~�@������CE�*�����YSOy���5��N<����E�q�7�y-�@_��-)���xꁉa�3���3]~O>ɎhSYa���wS$���LU��,*�	����B|�y^a����O���l�W]B��ț�o���}X>��Q"R�?��a��H�s�|�D����K !��ֵ��b����M�|�A)�
��ng�+���%������SM�?� fxt]6��(B/���N\li8� �y���ːUwa�ˊۚƨ����,�.�N6���K'&%���=��e���l���?���J��a'�fD�,��qOt?��z���8W33��-��gq=r�P�����)�d��#^2��|����K�fr��`��8 k��S��}�F�-��aI,�5����H)�A��?�6����}tgSe��1�.!����t�a������`+b�Y�2���O��� F���������7�?GG����^�es1~y2UM��a-Ґ'%CKX����V�N���K�Bnei��&@*"�^=��ƯO~y�)����P<��p@��#�
(+b>�$U���Ӭ!Yc#8�!�YwDv?F