XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?��ݩ�b"�(�M捻���,S�A��pJ�#�A��{��|��tT��J�Z�֝�6,]�^��`��ְ.�1cy�;Zin1 Z�x��7��M{��g��T�6N.�0ZALUlґ)�Bk.�Cz��R+��7[�z�I[Ȭi=l�
{�d&�#G� ���<ᢍӄ!7�V��(T0�����P>,:�c�Z( %C�y�n+�-y����[��=�[�)d<��u�ɂ�Oț�W����[J b>���.E�h7���D�AY*_��D�\���A��éI��r��r�Yv�	�U�p�J��<��  W=�����!�m�#��-����$��pi����'ॵP���4e���~Ĝ�Z�8�t�"���Ke�t�!Ԭ�.{�2a�)�lA�&�Y���lG-87}��f�l��}�pWص�����f�[�f�1!y����q����7��\�*a9a��r 㔺ywÛ���T���E�!�d���@�,2�\B��rT5o�6ʹ��h7�'�Dc��Bߎl�[\1[��5B^�F�H�����ϸb�Mk��J9ᖗ��%�Ick��J:�{�ҏލ�+����(�<J���˻#zE]lȉ>?Sl��]X�\�ne��5;��`>fR��[���a��s��x)9_�� o|8��X�,�lJ&�#�2�G�*.��s�MY����*�y��	m	�D���q`d�q�Z�f�l�!�P��p�N�A��˜ۜ�9�})�����cp�%�Ӣ��aIgUQ-XlxVHYEB    3a15     d40ܦ���WC��rhup�}�Fe�o�b��7�1����I=&v�K�O�,�(9d�:3L�����Fy���+G�4Aֵ�jK�B��px+��S����'�v*N����i� �4��H����oA� M�vp�+���/#�%�U�j�N�V��C��,@����RPB3&����m��.72���wJ���Q�H��w�DV���� �Ӱ�k����AK|��Ӹ�tf�l��Lc��B��Յ�d�3��8��>�%�;�l��h}�ǭY�J�����tX�g�Iy��� B���`�"�"B|��;��H��ʕ�1 %�U^��{��OrDi�_8;�����Wi� �$�gOQ�&ߘ�uXo2!9�)i
�}"�]��2��"�mu'�Y0]���^,�����@f�vۥP�d�o?�W��k;�L�B�7x�i�:�^-��6=�5G��x���M>�K�u�@���;v�&�%&�;��{���q'�}���;	e&�\hd�(-m��F��Kum�w�tM\(K�C=��¬9꣞"��m�lbK��!AW�k�R�l�F���L��m��$�R�`9���ѣY;�&[���y�C���+-�eH���G�t��E�� *P������8}X���Y���
�<ڌ,.�֎ZƬ��P��B���Qi�.��n�B��_�["��]�W��2��v�����-ݬ��=K̀CN��� 5�M��4P�_}.	͊�`�����9�e����s�#O�yIYՂ�����l�$g/XΎ�͕k[�1$�f�.��b����D�-WyŠ�v���Ge����eZ���+-��I�v����484�D��?���b��S���\��L<b�M\�Ñ�J��2~�3�8�p:�o6�\f�;���3�Q�]��~�ċ���atBJ��a����U|������ M%8�@�b~Ļ,ı�D0wR6ɟ����1����y����,��/a�r��?"�/�b�V,$d6��s��
Y�*	�-�����.��c�ɼ�n�Qt�R�v�T�)f724E0:F`�z�����N�HB��O5*
�%��Nڀd�.-pH�F8���,�����$���(s�t��LU2���+j�\%qﴼS^����v7��^�(���LiW�6�/���b̤G�7c�FY%Ľ���Z��@��7����i?�F�����o|"�W��x��[qm͌��|s�c�L�S$S�Tvy��[W'�h��dz�[v��W�4��{�]10d��_%7��-���4�jr�%%�[���pҕ`m=�	��}6�ߺ���I�c��4qS���;�ZۭT?�&�Ay|ڇ*�H�r�#��O^��).(�.�2��wd��m��\�$��a+��(�
�]��j�<	}.��i�����عi��������S;�澤?]���|!� ��f�
y�7X��WKx���"I&M~��z��i ���_��;;RiI����E�&?ʹ���������5��mJӇ:�op����[��V��l�!��O�����/�?=���<r~v��U���@q��y��U֙:�+�H>p�o
���ʹ��Pz.m>�x"T��6�_}�W�ww�����:!���o*���Ʃ�W�!ڳ�V�_O�s�z�걚ݢ,�i�f�T�,������Ԡ�A�.�"Ab�*�?�(Wf�CzE��K��CE��������A�#��?���B��Wp�qY���.�a�R֞�Da������D~��:����!q����BUj�y#��م=���\�JC�O���yV�3�/<�-����/�6�*c4m��d���x괚�7W�pH}�M\,�u9O�1�&P��C�jĕv3�D��e]	3��Z���?^I��T�$�*l�@;�Dr�������b�+6:5�xDq� ��BG�C;�'k6/��@	�p�{w��z�`v�5v���2�s��u�d�p��3�'��\��b�L�.�(���2������RHt9[�0�EN���~"���刲3��O�����F���RX��[�w�m^6H��]-�o��A�}~z�&�#��̊L;����юSG���O�T4DV�6��TPl�q�a)א�k`����f��4
Qv������W�+f\\��޲O��N%e���`G̡�J�aӫ7�{��dSRxT�]�Úm@ܽ�+zq�h�KD0���ɬF4T�K����2�����ߝ��hf6��9c��Tiy	l:�x�C\�l$�jb���	}��,�-�~"п�T:qM�>�˥^�� �p6k#.t%G���B�{VIuF$�=V����u�;k����DC�G���Z܀	���\��em�&��.��,���z$'$����v!���H9�3s.+׿����{
�z����lF����bP������a���1�ɮ|�h�ӏ��wocA?����?���,�pP��)�@���8#��ҿ��(t׬�STу�\�\a�!�n�����V�>�H}"�1�"�#�Pf9Am<��n��XR�(�{�'p����غ&̉	�y5�O>H0�g�s۴��v�}����-��7>����+��>���~�=Q�D�Ͷ����c
�[SθgN�حA f]�1^��^9'�tM��c ��}�^����*���?C��̠���y�������E�h2Y�EJ&h��j���w5��!�`��q����G��*i�fp�B����/�W��pɮ�Y@�X<R��YEty�R��9��׷�ДbC{nLÉ��[��Ԭ���@y`h�$iH6O�)f�/Xg�~pH	�I0S4�w	�-���oc���迲7Z&/��!��F��6���Ot*Xx��ů{V�����)Z�r�����ym)(;��5$���M�?Ne��A~�[�l��7̣�V�CK�
_;	�m���Ư	ﶙm�I"
�>Թ�ㄓC\&�iX��C�~���S����7�T'���v�.�(u��d�Q� �	��Zp�ZǛ�8�*��NL��� ��T~5�4G;��N�
<)S��|�O^��6���s�Ѡ�4��ʽ�[��7t�����?(�a�ar���а}��kkXq���!�="˔aG�]óʒ^;<�w����Ƥ�m͏EK-s\�)� 0:��9|Q�7�+��ƈ:H��L��̪ܸ�p�X�>�-ר�^-a��h~�K���F�wZ^���X�n�s��3��JqKy��o76�@����@����@��ǁ��˪�5ޕ/�(P����ۼ;�+���?#v���e�e�p����x=⥞��Z>*�p��{`2V�C��Ģ��̔��<