XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G�Q)Uېj�-�z(@{2�}+�#���H�OF�A�$�"[�Ƭ�Ҷ��4V��?:iH��l~L7N���Cl�Ɛ�b8�<�H���L����l���R���C4ȸ�d�M�v��L'vVy,&C�)q��j43c��3ʧ%�tic�aę�01CIfgX�]d,K��C>��wgWS�������o���jof�
%&s='BF|(���e&>K����B��_!>�]1�;M����@"��uy�%���+�
��{�z�{9|�B��Q]�<�;p����F��0���Gn5[%m�MLZSN!��bq�l<���JF1������Bp��O��-���OkM�z���h�SĎƽ|9�/fD�4b|bT�Hu��7g�J����"�Bf���6<�=�]��(�$����Q�ݠ��~���aP��{��+���g3�}��P�ϲ�}ndi��Aa`C�[)��L�J����Pn~\9�,9~��s�W�Ǡ$�<��aHg.������Ɏ���j�j;-Kc�4��b�1%��"�>��3H��a�u'�t��u�Z�|�W>�6ϨA,��(g��Ra�����̲�T��R.4�,�%m�Ia��C��?[�5	�H#�unnn#\�е���f&�{U��{gy�r;��������zx�1?���x��pL��ZNG6 #~9��]���H-��Z;zm~jy%Lެ5P	E��gs�V"jk_,/�AX��X�-05

�A�����"K���ɅXlxVHYEB     6ee     2e0�(���i|K:�͞|���-�Խ1�0�dh%r:(�n8Ǚ&�^�(����G��n
�SC��=Zo���B�q�G�l�2�9�6�5��H2J���Z��u}=It��w��	d�2ȷ�$dP9��QM����=�@��w�^���n�����R/���?f����
�δp)|���a`��l�YǨ�/�(���%уo��E�,��N�n���^y����s%K�a���zM�q;
M��/��O`�ջ�/%Y���t��o^�~tHV����
�f��a~�\��r����bb�XJ	Z��?��sw��"�	�vh��I�L����e&��ǐ���4�x^R��Q�>��h��2<)5
9�G�n����'<��<E� �T�S�A>(��;�:}h���5��f.0+{l�&�ʸ"�CrEi����F��8!�u�"�%��[�̎
ĭ*[�^Z��w4��&�ƻ����Z�'�/JG���\��
�d����ʕ���65�v��<K >X�!��v�@rx>�{�"����'��D�?��t'���a�l@88�xdwh.*�o���R�P�H�yn���(�Ž\q揋:&1��f�>��C����ҠA�+�Q��.pa���\���;u�I��C��!2��w�,#+o?$�����3+gk��[w��3�F��AGZr�8U1A&�9����pZ7�54�- ��,x���	Z�k��)VwR�