XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����BV�Ȗ�� !�Y��r�Ѵ�U���(�
0�k�?���ǁ[XNLl&4�È�N}�l�1"��=�e���y�ėш�ĕi�u)�N���(����HGl��{�u�OP`L�<J����y�x��6s_f�\�尰��^�%ct��\M��G,Kt_n��{�x�K�V%�?�S����7��y�=�\6���c5R==M����ЛM
�@�����,��b�����/����j���o��m�p ��fR:�����o.({�Eī��tU��d���]��h)��"�7�Y}!���-����S��D�@}�{0�t�4���6:���c�f��H맆/0�?�կdjN�P ������o���O~��*�Jb��-5�X�a�*��=�� ��|�@p9�BL@o�_R�t�Y �̡,�D�K��n�]ꏲf�/Ka�d�y3�Vk���r�D&�#!�XCG\�4��$���הP��IY�_jFa>��ɤ.�Ʒ��AYT�����wEʟ�ڴ��f�D"����f� �Ln�aq�����_.pV��u�j��}��������o���"CVuM���?|8A�d���QRdͪhƪ�f$YP[}�P�H�[������>��S�67�Wh��nܿ?�Y��}6a���=�����^�,�:��kS��G����@P}����ݹn�I�7���1�45w��������.�u����U1oҖ���	�2����=�2y$���e�YˬX9XlxVHYEB    165c     400!�D�����
�x�3)�Q�i�<0�!u�So�����Ĳ�m[3nN�^��@�<�SE%v��{Α턍��ǞK0����G��WD%�UN���+�4.��b$^���i�'i�UW����Tx� ��]� �3[���b|�	��g����K5x�}�&َ�ф/���zwM�ap�)S{}�2�B_�70>���n��(�'-G��'x�%�<5c���sD7����ea�%�����@K����kkz	s4jB��ˣ��$uUb�Op2m8O���:B��<?��'x'�����=��� "�f0����e�ŧb]�l���G�K��4r����$�&/�����h��r#&�x��,�I溇G='Y���u�Ė�Β�;�AL��*�l�Ч7�d�2�6�'*Ɯ"$�P��ĉ�=܊���9td�9�G�=}�I��\cڦh��Z�����0r�=4��Q�Ntw�����2o���b/���F ��SՓz��Z���R�\��(x��x��~��:4v'��� �1��w�g�牼��*��,V�,��C�G�
2ㄣx�c7��f�S�A���XZd����Ms7�Q�!9�������$9#�'I�pmx�H#ʾ�7��RZ�u4��!�5����<��Y�q��0퀚��o�l��5��v�7���0=��bF�s�qǆR�U����9�M�]�	���܍B-N��܄��
��6Z�`��^���*�tg�� Dg��_��!�����K��Sܙ{R}�%ֶ��ֶ��e1F�������YEP�ѣ�/A�Iжg�7���n=1Z�����M4Y��B��z�c+4���$fÈ�)!�o���l��GJ��r�2a�c~�CE�2���>�(#�`B���8�c�B4j~}��)�Kﱻ�l�{`%�[!wU۸7��.�1Ai?��GD�v݆�� ��)a}Ne?�QV��* 6�d�����b��6�]¨���H6+��0�t��.0-��p1��BU