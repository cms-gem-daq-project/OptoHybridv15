XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+��a�;�+Z�b�g8���Kk��ژ�Q��H^��`����y���Y�|�E�J@��.F���vW�&1��pd�PV�������6�i��E��)3p�	��WI���:@��_��m��ys�*z�"o��Jr����"p����?�u!K�?m�s<0\�GSV��9*W��"�v'��9u]��>쵻 �b<t�h��g���p�X2�D�8]�u��+�R�uh��I`q��ҏ�2Th٬ŅD��c��F'W�T��њ�#O�*ݷK�ܜ��C��¨�����HbR6��Ш0U{A:�`n�#1�*���3�K⏛�Cz$���ƚBͻ�X�	�v=�;
��`h�TU���d�-�m%��vKI�9V�~#���S�P|(��?��$���.[�GX����1,M$]���g�pOK�V3�kY2R]��#V�D���Qn�ѽ7B��$�iw\23����`K6�Z��^=�wY]KZ�,��]ZT�� qK}a�]�r���^p�`[Yf�V��������WE�?n�gZ?7�-(�n�)�{D��M�
����"G����B�I0��cO�|/���(3�Ќ����+>�ޕ�b򟪬��L�яeu$�̑��MS�I�N$�=ߥ�d���)Nڵ]ct �&�Ş97^��_���:���%���?�<�_�?Dv�X�Kd7}k��5i�v��#�3z��bO�h-�N��Y���;��6�<���f�t��z��K��˘XlxVHYEB     6c5     300��`r���ٺ?v�'L\v�hy�a�r�ͷ��R�<㭉�:Xq����l���C?��AY`���b�rX���v81t�o�u]p{���?�A�������v������ ���˨���<��g�� 6�#s�BF�O�>?�6�g��s��0�����N:0���۞������m�2�K�2`�vUd��3��D��D�v-�,��n�����L���]�6������0�J�a����vk�7���X��z�G�M�7~�2�Qw�
��*�j�0C���R�.\ёw;`����,��O@��؈��s,"����KB���,NEt�Ό?�p�R��)8�2�L��̐���:	�V�t՛���C,�٢P�iF�p��d�nF�m�xJ�F��"P>��t?2w�O���P���������p���rfΰ��k��m)����R�����~�Ф30�l�Ù\�G!m���@�� d^�>\��"v��S8�[í�D��h.���.��L��El}±��s�c�M���ZU'�r��(��pTZ����F�+w�k��C���v �#"[}sx��cZ�}<s���mr��V�T�|� 7ʳ7�:2�
uCڐ'�{���?5���Sw4#UO���]��Պ·Zs�M��+�)���FBc�{����`N��=�����u$(�_�@
���P:oC-F���������� ��~oí��`;�{LA�e�V�o��IZ*QcÓ� 	