XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��SR�����c|
����<��i3�wp���� �	:aH�U#ά�� 	; _!��������^������D%<�UU��!Ba�b=�7s�R��&�"�b������Bw�:��M���[�|�]�����K+k���1�����q�5��X�++hH����W�\&�9J <~���F��m��g�jU�G��Dgd�{[�#�7Q�`�E�T?�Qd��յq�O�i�w�����fx��݌x��CTl]��/{Z��t83����J�W� g�$O�m��Uؔ}���
�̕LyG�&D�m� �-��!�%��t�`9]OB����-�KeF
@��9�9�U���O]��E?
�?�������8 �ݽx�*��\�O���y��Ed�ޔ ؏��@B?��4=	������}����2$��7=ns�����a��Ax�f{NbF�v�������fT�-�H��|i�U�ˡ�\�����!��.�j,&�c͗�{��-�b}7�[��"��4�K2���F|�=1�@o]H�z��dϟ<�b>xA��a��J0E�I!k�'��c sx�^��L#J[m�,��;�eν�R^��ȡ�3�&�'�v����]v��:tƸ^�}�11!9[/��¹��X4�AǼ��_k��FPzr̷c�L��x�^Q�:Qk������#�V�$p�c�I������F�}z�x��E��<�f+edw��/�Ѿ��� ��G�t���
�+��XlxVHYEB    41cf     c40Ys��i��鐱��<�=�y�/B#���tD���DZ�%G�P��������B�Kx �&����XΚܢ�NE�Y����+�����D�	eu��:�'�rz�tѯ��Ի�n�s3��+�W�^'d��~��
�'7�;\����Q���b*���k*�;��묁�Hs��,�xx��WO>چ�5!��c��� )��x;�����3P�\Ѱ�g�M�k(]�!]y�k��u��\j��R��ɥ{�\}(�:c4ݮ�ɂ����6i��%�-~��0���J�� �(j[D9<1U�|�)eG��O���W�z���0��8�Jy�f�Q��Q��ѐiұ�n�NзE^����)<9.T�8��'O�&�
'O��9�N�������cE�|��Il����<C%�VlO�廂�?��^����Gx]����͉�K�pXyp(#$D4k~�/���m9a�3���������;��m�  ��h#���MP�֗;���7�&�Wx���d�PR�k,-�c	П�g�����R�4���֛����;a���z����.$>Ea��q��b"����r�,�����`��O�X0c����幥 ��Sy���x\P�,Gx����86?�ܓ��Xg�Pau�6��Y����0.dP,F�	e!+L�(��$1���PD\W�H+���Ί�+Œ�1��O;Z�i(n�Ħ�;j�tr� ����Z��������R����ko�7�L��������ѥ��ka��; �k�s�o5���Fd�"(AnY�1`!7��`%�m�o:�#.Ӆ(�2� Px��;cjz��z�&��A�l+E[�Y<�^��t�AY�]���'�⊅1L�]нK�]LA������.���kr��;�^4��Y�(�ys�O�O���hb4�\������(����Q��y�� �7d�?�a}����)I�0��s���:�4s�<U @	�Zdd�Q�,� ����揪?�̥���X�-*�Oxl/y�a��"��(7`��05��l*�ю���׌ 0���&�#��ފ�|�-�J��mM�0ϧ��\����������O�/��J
�^Yڊn�ߘ~Uh:�$������-?eԢp�ڋ�� �46z�&�J������в�eO��>�v�ܰ�6�#m�q�,�ef�{7b��d�~%yX�����OE��0�O��2��'4��@���!-YO�F�}��/"j;ק'*�m�9�f��n�PF��C�6����掗x���'F�2V��6�n�w�\�d�����7�����Bլ�3gR�*�2j����`�.�Ǟf=�>3�"�
�~����h4��)�*\t�+{��0�]a�����3��Ò��ƻah�~]�l�bY�x�����PrB��Z�Ww�!i�O+�-B8�Ѓ�v D��aj�O��<�}]ߨ�2����d���5�s�ڵ��9�?56VE�����O�ߤ�[��Y`��q�¤��b3{�m���vHfS���ٿ�#j;$�D@��#񙘢�����zUdn��޲�u
@�|����v:p,�6;gU��u���%��u�a��d��t-��V^{Y`Y+:�����R�����Y�����iu�7�������bU�CEw�ֶ�0'H�}]�O8I�3���K���U5!�,���k9��k`h���de�Rz����qT��eE�J<b1'���0H�B��bZ��-0��\�ǁ а��D�<����Qw�.���49P̽�x�� \⧂yN�hz
^�'=�4���/B�O�ɖ'.��FCt�ԩ��$H\is�-W1��ۉ�lSe4^���󭂧J�@���׽�H�_��z�+����]�׋&��,@��Edǻ���e�ꛃ���O���w�bv�zb)BL+āt�A*��J�ǘ��k��� ��Y��(�]�*�c����T�� ���n.�������?�P!��kxN����숿&�� ����-ؓ�(ɘ{��9�#>$�j�`�W���y�Jjȡ�o�U��³j�*�ȩ7�ػ��iKW7w)T���m��)�,og�:l�)���>����a��pl8�Wf�hkM)�ۺ!�G�o���G$:�7��jԜ��.����"� �3E#��� rP�ƫtL�My� U �7QXO[
9R�E2jV�J��l��͑�n�U�L�K�h7�63��J�CH��:��!��_�'ǌ n�*�W i�h-�=}2JX��-Q���`A����)	7�*�p�Z�r��2�8Huf'.B�*�?����)���{�T�H�TǠv�?��=Wze��_W��yH�F�)^�8�y��R�[�(r���K���#��-%�9-w����O���1�Q���>^��3��fc[���={���%�-�<U	a�7��1��/D� y��{���H���dA�����B9ʅW����r}�LH�ҏmr$�`|��T���2vb��
)3��<c�q�������'��;�Q�NZ1]2K��-ޛxbb|��;Q&�:�b�h&jR/�cC����A���K��@{7�c���3���/acF�N�E�o���m�l��?٨-�<^��n|*�y`J"����C�1�B����k���aQs�.1Z"2���|�Y/���1�&�Ղ�9��7X�� ���a���a�ǡ�`/���IժZD��G��>{CF�U�4���XLQ*}�x�\Ǧ�Г_�LY��R�I!�Ɵm/�k���R�[�1�O)#��jPJ������f�����T�Y
}_�n�o4�BӉx�/�G��}x���
ߜ*�0؆��cA�_�l����E���:<�#Mpyu)WAB�L���r�I>%�C�pl\$���U��7=]�� <�M��9c���6�u�:F=loq�0?������K@pL��/؄�*nB��
�-R� �o���եAAHeS�q��(nPT��*�Q�ŷ0.�*f��&,�S!a^��8����]ĳ�"��� ���%¤*�L	��=D�f�p:Ah�4�B�	/��w	��>�λ\��$���O�ꬬ9�*���4�,�=7�8rg�*YhD�O�