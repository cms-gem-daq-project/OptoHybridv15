XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W>4�Ψ��&ڶt�<'�U�J�LB��S���ҥq���]�RC�ƣͿY�&p��<���_�}q�R���<�IUǹJl��ς�ƾI�h���H��ϓ���ǟ���:� 	��;�`�F$OY����fL$]:]k�Y6��~F�p�+�\3;i�SO񑸯��+'ޤ�?ib���w:��bH��3Q��1#̵Y���S&�d�(B�C�"�y.������q��3	^�����/�ɵ�.
۱�r?-U9��T%��oV�rʙW��c`�x�3�ⵞ��"��lC2��YzkƋ��SQ�/�M��l�>x��YF��G�M��׵���Eo�]0QtUM���x��~[a�)��R�O���<�\�=r�5a��{x�h��	��c�?rr!F�Q�[��1Rc}-	1�0m��q�賾_Г�|Ct#WDY��P�sEt��+�d|�G�����%�|���o���J��jOq����k%�)6�ȼ���"�߳�j�3x���RՁD�U�S*[~�y_�[��?~�3N0}��p8|@���y��pK#��.��=���X@��Izr2w:O����ȇO���!��۾��988"#��J�e�y`dp�j�2�gG/���M�ڶ��9�n[�LM�#z`hT~lQі���j#Mf|���ep��w3`Β-� �2��oc�c��� 8���-L��t� �\^P�T��������P.>nwq�U�E�L��[���\>>�����NU�AXlxVHYEB     82a     300}�@����0�z��c7�`V��/4�'�ۄ��7��ț��Ge؊cTS.>���UpƲj�sE3���0@�C��`���-;��R�]	�C[f(�¼�57�3y=^��,x|݊�Ϩ��n^Fб-�a�˗x�=�h)�	C���D�I�l|
���8��2���(Og������TL灭�+o���'Xs�$0���v�6PԸ�Uh_^�]���h�Pn�+��W7�(C��5��s&�($L_� �O���)>4����i��[Cy�[�C�e�uN��KYd�a��=�V(/V�����d�H�$�"�-:�<��nʬ�Y&M��-W���XuN�=���p>�iFh0�����]�7��;��A$s�1.}��{�[�6/t��~���>��5qh\x{Z�>q���A��1�W1��7.V+B�,�U	q�iGa[nȔ҂>~��6exn�yP?� P��j,� ��Y��5��l�*�!S�ɳ}̧�\����bչ8����H�F����'����s�;c������w#\��?|n8ޡC��@���'��EƄ��F��ˊ�=U79���[��ń{F�;+��EW�7���]hO��� ))b���'b�v�oWՉ����k�����k�?��xS�,odTn�l��<�棑�(��~+(��;�3��T���l����+�u`�����:+��h����V_`��>ڕWʿx�d�1Rr��R�ԇ*�y��2Y��3�u�Fy��m�^���g