XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���BN7��YW�)��5-��q3ߞ��_Xp?~��ÉC���"�L��7�5@ t٨�+�n����c>̏^8 �6Ѹ'(�v��j䛡�P���u�W�#��O琯���q!��������K_,��e�W"Jg�3{�5�!�g&p�c�FҴ����� ��zsP�e�5��������^�֩�T8�q�w/A)e��QFԍa�c홣��i�׉%]�#%�v��L��\mWjI�eE5}�=^|��D�ǉ��Ao9��Q�J�;��]�F�89j��`!�5'h�I��5_s 3���V�a��t(�yJ���&4���t��d��oFջ�f|����GgFR��zzi,!dy��=�2�B#D@'MO��'��VT}��b>�~��4��ͱ Y�����u�Jr�UڽA�p[y���k�"��qT���9э�BOFY����L��c�Q����1�(Q��I�>p�[���p�R�T��g�G�pW Z����H?R���ƺ�̍���N��� u���t�_'�l���4\�EZ�[��V��-�Ԛ��:���RΞ�VK��KǛ��#a�S��YQ�C�֠�ۜ�~l:02�B���:��*|����������.���\C�,p���'_��E�٫��(^(��a�`{67�a��4����2�C�4�a�u�-�8���SsX^�c�L�_)�XjЮ�T��&oM	�L�b�3qO'9�Z7����Xni;��[����T�� �w��^$|�鄊s�SXlxVHYEB     d49     3b0n�~�	��Ne�������
X/��T<��'�~�À$=�ړ��+[��A#�&̝$�G,��D�}҄�K"����1�����y����8��]� ���:��Z�ew}ۢMVSE������l�J4���Y������q�����`:J�p�UZ�8�o� �U�אu6i�n��,����N($�c�.M�i$y��#ل��DF����a�ȗ�̓�/��)�-�:�)`��RX� ��(	���b
�5ߦ�>ߨ�٭>R�{�	�4b�t��{�y
�7��a5�w�_"�$eD���`�d(����X)����q%�ؐ7ۻ�Oj^|'I+͡�S�>$u�Aʺ!���� Ǯв��莑̮�\%:kV~�v�}i�/�!|#%D�q�R��ɻ<�ihoF�n
�Q�#��T�;��n(dڥ.�[)x�Y\�g��f�Jf�Dӗ3>�_m��#1<
HhY�:_)�>���-�Z2 2����w6���]�H��)Ҟv�p\�Jr�P2f ���wh�+�c�yFNkg� ֫H.[������'���z9k�_$�(�+�v�vc�\K��܉�R�n�^rZ87�'��'\��waV�R���PccH�:��M�]Uk���u�c@�fZuQ��)h�e���o���`��l a�X��?����,)!�?V���,V��	y{�$�p%��W�%���<3�&Y��l�GmY-O?(X15/;)ɞN,.��J�Q(��kF�D�ʎ�^+~�2�ݸ�m��Cs� /R�'Z"�a� �;F�����R��,�A���9�zt�h�����n�|��DFN!匌5��4��z���Rn����i���&eD��Y�hU_�Ǯk\E�x�~"|�U�rh�O۷�S���gBS��L��xI��y��銏\�eH����PۄQ��=�W�ҘK��=Y�BJX8.