XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.���|�=Aތ`jg1��O��+����R�o}	����8���屮�l�V�$c�c�ǣP
ez�-��f�s��?�Hcu������:��	h:'^��.$T�u�m$�я>"]�3k�9�h��������}��03@1�5�:=�I��<�P�Ш�� ��!�يʠo�I����7�fAFwh�D}��sܒ�������,�L�A���w����\�R�y�\�	��A�蠬�B�}̦1��N�f��l�E�2��em�9���T�u���V���Q����8
�x�p��Ƒs0=��KX���r�DI9�A�)�olj���B�̪��@�l�1)Yڏ�������o�gx����^�0��'��qQ�	�yMr�	S�k"����WZ�1'6޸��HHvI)G]	��^�:8�Tf1�Y ��O۾�zaʴ��|��b}>�����R� ލ��3��������@���ΡT�$wJ���HlQ��{��}��w0���rB4p�q����SꈮV��ϩto���I���mÒz��W�<~��k<�%`��c�'+��_MtI;�es��G��+���/dfW�0 ����`k)Z���M��%:,,��|->��w.lNuʙ 8SM18����R��q�}B�G�����V�Ie^ �̉j�0� Q��{Wf`��(�S���cH�Bt�O�Vg>�E����qCy{<|fH���{+B<-kb���M'�/�7��n62 k�1���2Pd	�XlxVHYEB     9cb     230`����Y�[o1T����o�ۉgq���k���̨Kb!�����.��zd옡���1��	��u�*d��P���Ux�oR���<���`�D�V��d���1I�q�����Ui�+м��WK�@5s�
#I.H[�ì�K�Fa������-ˬ8(H�,��kqq�Ë���ƥ汲�����!F��9�Y�a�����ڭ�����e ��Y��u���{�܃�@�Cj�ou��<E
m"�Bf`T�7Q��#s?��ʹ��}}	qTfI���̥+�ީ��Oso���+�5I�䇯�w�lp�A�Yw�	�>1\<�C�J fdy?�v�"s�~,-�ڹ����|����S#r�r��F�F�F �B�(��r�P��jv�Q�I\�8���b�����I�����o�e
�w�i�gg
�W0u��=�`ҙm��[G�+%�Q'V{�M������.䏴�He��	�w��a�X=�v�� �`����c��^�����I��XT[l����#`b�x.s��q��P���vtظm��3