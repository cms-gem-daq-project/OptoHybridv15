XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(����0��rj))�|�J�[O�7d����/� ?�z�Ԁ�՛����`^����dC5��K��D��( و5���K����e�'TD`��N�h"�Y<v��σ݂\�f����M2�U"���$�@�DK}�GDE�;��]b?*�z�&��I"���?m�]�'V[}��cFXQ����ȓ���pO
'=��6�xO�?ȫ��Mm�͋�A�6�	m�I�w���q@ֽFo�Hf�������.�c�L����䵶 ��,�sg�!y�u��%R��Z

��Ҋ���x+�j�ݤ���[��R�9�J��W�h�c�t�dB����8\�n�؂�����J�69�p֨�`8���6pg�&�|�
�����U��bP����׀t���mQ���|�h�15Q���0 N���tc�d�NT��N�6�0a�8\Pm��቗���\�w�>{ɕ�$؃u�}����A���m>�ڗ0��c�i��[!��j�(������>�sm,� E��MlWh����iߩPS-���"���~b����*�F�?��.��g��]�����g���z7R/G1�������kw��)�/�ggs�օm�@9w)��*�|=N'!�@T�������j��CW;C��$}��������ǿ�ĿA�f!�[��S�K�jR�	M4���Hn(vuj��=I��7b�3�0�v��Yl��aL�-}�3���Cv��fJI�S*�I�]k &�e<?:F���ߍ;�ԠSKލbX!?XlxVHYEB    6408     e20����$������9������w�Qx�"'T��q5r��Rto�l���D�sxt��0Ӏ�F.�u���ϘJ���.���s��9�
\�ʭ���]@��.��'�E��Z�#C�`\_kdt)ou��i�(Δ���F��t�?�%�|k���tS��k��b���(�M�P�*��)��#����?E¤_l,���Tz��=���ļ>�DH��㍗��vvΪf�Qś^����,D�}�)�����'�2=#a��kgq�V2�wGc�+SN)����^�[^����eB
ŲV��g�o���~����^��D���� ���=V�2�j <r��1g��-z�����E��`,B�̰��"�m�W8�:p��߮ �3��],Z ɨ�oO�]J5i&RG�P֯v�wd�L��<�m`�B�	��}Hp��|ٴ֤��,�k���n���6�ǚ�qW��{�j�D���ʻ���1��(�o�~�88c7TY�R�A��X4)�մ/>�L\Ӂs{��ط?K��Fj^6�&�<d'�՜�H�\��X�繊_�j2�×��0��|����w=b"cp(��,L?��\ E�T���A�k� `/���;&?��[��o���d#�������＾�@��s����	���5��y[�����DA�����H��cc
M)*�c�/;}�DZ�!�7�y2h��,=����q['�ͫ�(�2�/o��@ư1�j���J̶�q���c3�(�3k����@� Eq<���8H`�="���<џ#�,�d����m`�6���z4�,�Z�p3Y��]�vgR����&�5J����Yt��L�1O)�^���=�Q��N��♓���G?$rf��F-u"��)J�3��ϒ?�*}��*Njf�����l�Ȇ�|#e�ll�z�}��rj���:�|�%�Ҕ3�Ot���Q$Ϳ�;Q��Ľ`ې@�Y�P���z��'�����7C�us�/�.uo�F�% pI:��̡��04����;k�2�4�P}�˕r��.zg����+-8`4�Jc��TDM̙����]�;�/9�E�-�U��c���7��ۭ���μ�pS�������^Ś���?cG;�u
V�LX�,C��
�w˃�v��d0�l0��fy�R�^���'4ƥ�}^�Yk����WsD�nx�9B(VҨKR-Ob���!��WrB[�5��nko��ی?�^Hne���0��:��67�ZI�(`,A��U�F�>�Vj��}�i��������7���þ|�	�_뻧Kt�\�7凜�����#���:���^��=�s��j3�/��"��Ŝ��T��׭����h8� �U��ЕN���t��qu�i0���(������xa�*�7Q�˅���x`�e:�^��л�N�1�N��t��NK���F��UN�x� �l�� `}����\R���$�?5�H�~|xIUQY���#�
H���_M?Z͝�5@%��/ծ'�`���bh?���u��)=[1�?�8����:����CD��I�,�Y{|\��@��4˯A��kj�l�H���Jxɘ
j�a�sb�[`�G~���\�@g��Ur|Kd�����p��S>�����BL(1�:�4�W���0�����G��LO]Y`N�Y�L�oLg�2�,�R��s��/r-f�v���B5jO8ޤu���D�܏V ����2��[���a��1�m7�Mպ*��Z��;�Y�s �<ra�dN�����Ygy�+P�Ej�z��46#m�L0�+��-�3@�`&�Q�%��Gc~�\쭿���CB�y~�F��UX���7=�����(��a���G��u#ee�D�5�O.���IG7�'f�<{Ş1����G�`��Ra~b☺��ƕ�;��c�bP=���%vZ���~��:�|X�.���M`�UWI��%��P݀�2s>�
w'\�l>E|�Y?������x����+�=��W�yTu�7�\3c�� _#]9i֢����$v�4�n\>��[�<S�4�Ƙ�/g.ky5i*�h{l�c�+ �e�I$ B} u+M$��L-�K| `��c3��M"���|D���}Խ���0�h�Z����W�̓Z��9P��d�y4{݆c���O�(�����ep�d����ݟqJJ �h�O���K�\ݖ@����!�PlW9��T�+�"�ʪ>M9�ـY����@(�\ϳZ����vy���O~ܰ�m��{�>l�>@�nXJ�y9=*��B��q�a��|�Y��H�$:S�%wВ�T�k��^ S��X#��p�df��n�1Z5����Y�R~����n�"ٳT�PL��{���|�w��f́6
%s�'r��ZU dUz�AEU ���0����ˎ���]��x"1]��pۢ�fMW�g&���2A���0Q��OH��ˑ�����ǀ��x��e�&��:9�@����nx�����,*G�^k��AiJ�o����V�ê�����x9 �Tbz�2��4Z�E���<��O��2��-.�lu�� Wި�6����W��������'M,���9�ٶ��^l�C�,6�쾆�=�H��UXq����5b���.�ݹ��}F9�@i�J���sf\G[i� ʕ⦡|����v� %�����������(�D����G�0��l��|CTo�v�t=}٘����`W����,3DOJX��~8�[�NO��j�8�d�^h��
����iZA�dK�Y{@�������C~q.�7��+\=�SS�7m��bN�)���p�� �K2�+*�A�_�b��Y��T�Nف����r'�����k�8}�1ܪ��۠�s���,/�<������ʂ���V�����g�ĝI	_��`jsV G��X Q�m�~����h>u��	���'�[[BË�-����x��Q�Çc7�����X]�$M>t��w�髍�UX�$���:��3��6�b�{�aU1�}$ꅦ�pNB�pN�+�-�ƟiN�h�bs�п����P�<c�J�x ^��wҼ���'ډM-��ȇ�GU�z�2�8���;���M�[+�QVڠ.&8���Q�J3O�&��!�.����y�j~�������T��ϱ��Y�"�m���!4׵%��|�E���0r� ��(1&�� ���#BɈ!�r�ң�r �b4��|�t٨���&������jL+ �6��V�MKo�ٿ�;e���|�5>����C�g��2'���� �����F6��B~u"��7k;v�''NY�P�W�:8L��)" �A��������|�Qػٍ�lr7bba'����2ݲ*
��`�(P����i�\,��z�9E~�
Js�Z|6~[���x��t����،�*�rdU�iq�B��Z���s�C������|2���$���PJQ��@贎�7#C���(@q�e���=��k���AO@**i��*�D�����������ј����'�
뜑`"v�x��L�x�j��/.4��/0�ujFr�C�,Y�:P����