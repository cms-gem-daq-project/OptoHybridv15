XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ß:��\�"c�e
��ٓJ~& �4�M�����4b�r��`Z���V�.��!�������D�!��5�؈堝���g��p�mEＲ�ݷ�f-8���FM(L�����}^ݢ�q±[P2����V�z�����R���K�6a���.�J�" ��͋o�o
�_Qjgu3gWy�W#��"-C)�MAD�ՌNZ(O����ZI�M4[G/�"A��1���= K��a���Qt�z��͖����/�W�+,A�;G�Z�k��@�S+Rר�9q,O��V�g��[xN5\����
��m�?����k��z�ۚ�� ߫��\�F���"���N(}�E�Lِ�K��CSU�u�6S+Њ��W�6f�IK|��M��  ���d-�3&�t�
Bt�Y��%����9KG��*9��tmX<N����"d�WЙ���Bj�iQ���0E�V���'�� �bI���P�����ݦ��Ёn�Mq���4D�����N{˖eM�2�p�o�B�3o�\�E��Ėb3	l�
#"�ٸݠ������@ �g $�ሬ7\�{暁�F�>e�̯�-G@[������v��:�d��Jl@"o�r=˔��G�]��=�r��.�4�����0�ڲ�t`?��wg�k/�Hg!�'��L�I,֋�"!�^�H5=�/�X�$2��F�@���J��h�?rª��� 'O���˂1��1K���K.*�R]�7F2{p�4�V8<@��{��lXlxVHYEB    60e7     cd0ؠ�?r]be���Nj���;��ϛP�U��^��8��	��|�
׼Uؙ1�N1��ܼ�G�+�TVeW�ի��Wܐ�
Q�h�(�,�R�q�q��3��F�Fͳ�]�|������O�Hq��]�������ޘ��CbI����hL��[$i�����x�5F�,S΍�Mu6	�A�'��zG�U.'yx'���RK��cwT#C��#2�[��'��R=��yeF6��7<�?�;�F�r���fw�׮�ͣ1��zǑ0�����T��\ayȢfC*���C���H���	yy5����3l�E�D)�B���n�q:{F�l���<���T����v/�K�Pl���/��*��~S�'�u䱙������������� �`�Ų\�z�v�9�N�_ߣx}|L�o<9Ä�7�^�>vl��}�[}8a��l��}о�}��b�b��o��]	��3U�Bp��e�nǜ���#,52�s8���޵ueɶ�#��l�=�G�Z�.��3/a�و�e ��,�(?�G�g��_7jN&Jg,�1���񬐸E 2���F�"�ڡ�"���,�@~+�����<6DB�n���}[]�T�07�����ļmM8&m�Xʐ3��*���������.iþ"=�C�A��F�G(��\�����T:����a^��5���1���e����{3�����S��*�=d܉8�+2��B���,�TcdQ�8[FSIF(������j�]���%!��q|8��&XyW�J�|k��ӆ�� � �Df{H\<�6�[堩b���豻T*Hh=��� )�I[��IY��Ch��e*�u��$��Y��-!h�)��2ɑ��ݴ7����ц�j���/W��@}M���-CJ[��-���5�Ċn�L�������j&P�J���)�*p�a���#e�`e�ebJs�D�_�Ueo��V����~��2I��07�8�w����C�݊?$h?~pS�D��k���*ض��Y�����";��I�H*��Hm�
�om�璛��v�U�����/^@�D��`}��C,�'q?y`��XV(q��'����mT�&<���r$���SR,W�Cs�͒�\,fV�k�	:� ��jb����I*3�|��;�v�p�u���=
ZI���,�@�+K�τv4��5�]�U�״�wFn��h ^¼��f[���Vb�B��3��J6/�
̷���,�o�T���o'"���s5냘tS�ՍN��)!�CX�52��K\�<��w�sH�zz�)gC��aR�#����>���^V^I�G�����x���V%���-?�5=�����<������<�5������)�9���-$驊���w2u-�	׎�څ�ϑ�a��RA��Q��W맍�t81��j!M�W�[a(fd��z���j�7,#-�/kW���Mv���1Y��~o�C��.nSҾ3�qV��:�Q�A�Ox��-�u��ׂ���I�cf*�xQL�Q̔>�)2�\�m^ѭ�=*<��C��Y^x=��Q%��v)2~�AI��GE;�S�\�E�2�Y�ɏ�`�4�o��8Ҽc5Z!�������*�hE��#S�u���BJ�l[�� �?=������"v��N���(�7Xͼ�<����惑�� Z<�L��S�/i̱4�����ߖt�Ǐ�8#�Q�:2�L��q�؏hK4�9���� ,C�
�b����:hH��U$?��l]6�h\��[�E��Rb�"�1��[�eߜ�;�[\~��g�M�gZt ��-	�^�l�YPf�_����JV\��
���]���ݺ��J�� ~2�.��l��h�}Y'T�2�j�����uW�����P�6o5�9p��Q�W��R��T/�N{�M�+��OmY�� �?/�&�Ď��&$bߓo��y؈��$=�(��;��U��7L�˄(/e\զ棳�$�v���v�C��4fw�i�A�tFM�f���L����xa����4�3�oಖ�F��g]=�U^�I�
 ���ΩՑ�rk��
 �i�M���1�7 ld���]G*� g�%F���}��<���Z�}Z[d�	,�����ua�<1�m��>tFֈ�Nf�}�� �?����#_��s�	GdyɅ�>f�Ncu�+6Ra>:
�Ƴe�91J&�W�}�r�u�������Ngp�7��T,M� :<g�E5��I Մ�bUQ�Cm66D�2U�՞���/�p�ޟT�i�G&����;���U�~N̠�^Ζ ���$%W?%6����U�%!�J���.F@��A=�v�--��(�}嶱��Ͷ�>jεx�󫏝�2��Uݨ+;m�%�P�1��9e�M�K�K���߃~��b˽�������aD$Sז�7�gfoK�Se4$�S}�ݱ�aY�>�-��VE�u����`D�h�Y/��w�gLԞ�Z�問	 0����%U�s���a�>5���¡�v�;_��A�hM*av��C��Ђ��f���z4�)�@5xJX/�=�PBP��){1%�θhd�	O`��B���E�a�s�l9�7NP�;�BMt�Vay����;�໙���ν���3���l!e���7ҽ��������<�)�:^�����?4D�%�8$������<������E���*���U���i6� ,�~����G��mq�h�F�yH�RK�9�<ρ��>��uܩ� �/�H�WSVGe '�A�T��r��1q�ȁ,��p�rj_��4hn�$i1%�{������@Д��7H�eԲ_�`�����\t�m�*}�㭏��cj�0�2GuR}���N2v�E�x����"��s^V&���:�״�XV� 8�o���2&��Nq�D��*�K�r�դPAW�
����uL{ג���*J�~{���̔���fE�*׊Nۊ�)]���ML���{��P�R�ceD c�5@q?H_N�P��S��]�����!��(Ƨ�'�����/&���Z.���U1ї_��ӎKfS΢E�_C�8L��f0sR��0������F%^���;Z�N�;����>��������)/�Ŵ��" �G\�:�nE7��4^NTo�6��.
c�qEz5T��h$������+� �|�.ps�qU����~3]���5�7����eb�]t�)|G��>��z@��h�d�>�d�v�?�p���$~;/��_�ٵ��K%�ە�yFu��iH