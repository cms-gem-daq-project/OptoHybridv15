XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/“��ۧE�Q���wɎW��8J��/o��C���:��]n
�8ґ����K{d��u�#��Q�$�e['���3�e7��jcHƧ��$�_Aa#3���P*|oG�y�o��%2��Zz�w��ٺ��	�Q$[���4B�(j�������aq|:uu
�a�V���.CN�ɶg)�k�K[Ԧ��̎�e��E��^=�&]���1��Q%���Z�H<7�M�Tԥ|r=�`�R�7�?0= �Uէ���5�s��Y�BH�L��
'q(?Ֆj�{&�5�By�����_�8�{P���{X�y��RL�!�gʥ���H|W�z\l�S���2�rN�K'bʏ~:�� ��R�N~�G����t�D���{��Z�'��I�~�ǧM:!���)K�%(O�y�7#�s�t��c�t��xVFb*�`��hї17$��i�ÛƼ@;�vl�7Z����4CǱL[�6�_��t^�&m h����!䷰֔s�[WGh���b\bEkT2��^V.t����Jޔ,��d]�ӵbg�!�%��]G )���ro���*���_F����坥���Df9Z_�A۫�OcY��N#@0��e���� Vz�/��'���F��>�� g������d���5bY�m�������xУsp}�KȒ��e-�ș��6�b�-�DK�[�[�h�:aI�2�Pw�y�&w��<��t<���POV)9�6陡N|_�$�?Uu��߳��KU6kֵ�=I��
���3@XlxVHYEB     748     310?��-�k�p��iQT)�A/�ZhR ��OyZ�ֳV-��6[g$��pV�����+�g��/���ڢ���������}��Hޫ��'����F��>v@�y�'�&����	YUt�N;���U�ь�nv�@@&ȅ҇����+�p���
�S%{Fȓ�j�0�w{8*�`��%� ���2����q�$��^�nH�{uϡFٟc���IX@)οa�uaOLdS��ˈ1�Nc�y�]F�T�F�y$�Y�A$���鑷���w�
���e����ܷY8m�@��P���h�%B��:�j9F0�R��������T��~��,�H$&��喜rxt�'G��� ��?�P�ڔG.-\�1!A���T�}���lO�q�d)����K,DB'6���̟��>�Ta��#��E�W}��ࡕm¶��!3�š�w��״
�h�E��.�����NB*E��h��a<k��[�3�<�	1���)x��na q�R}3��ѭ��L��[,��*�Eۡ�]-%~�3�Ս���b��)�d��}�ġɦ����W���K�l�q=t]Aǚ��TK�Ғe�1�~�Z�N�S?[���6�+L�nI�v8��p��5�ª�W-^����g��z�P*Q����ϔGZ�2��L��VL�������*2Z,u|�K��M��nL��n+»��T����a:�DpC��tdg�r��C�4�?caW�J���n�e�F�������h�������|۬���t�����