XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����"94�����Xx�E%�"�6b��%���_H��b��*xZ���A��'���B�Tu�؋&%`��8�Y}B��:v�Z
��e��X���F�A��|(�
\%7�c���!f���$l7Ll�r���-	��IpvMm��[`�GC�f;>4��P��\����4��ʾ�=g�șV�B`��C����0a
|k�A�v��m�����L�6x_.�&�qu��A�C)�3vň�/j_4�M~3����Cm_�"��q΅1��K��]�\�m�/��~\�*�d��9����$��,؍Ğ�_���5�k�Њ���p��?�r��p��'+�d��;e�E�7���<�X"�mX 泈��A8�W���_��������J�(����O�M긝d>�3��V�>�L4�i�m��=
��朅���$�Y]2�B˸��fT�֛�_��(4\T��$Q���.���8�5,���F���d�Z頋Z���[avo����eq�;����&�LpZ���8P�ԉs$z��H2��:Z?%g{'���Dk�=t��ם���;��̵.���c[h^�
�1H�re�|,fy��x:����������aڌU?���$����$�m���^����>2gʨ k�c�H��o����bר�`8z����ܪ�{+E�L�C��L�&p��:Ct?]�몔�#�����@J�1��[y��b��V�j׍dtHq~���x�������Ȫ��P�q�G��XlxVHYEB    b892    1b20�2s�1mALB��z�U	������Nb"�i����Έ(O���(O$o���h�^2�E1�t�9e�t8��l1[�A���:�ȡ�zI�d=�x���*�C�bMno����щ�aMIۺ�H������=\w �8 �>{�n˝IfX	k�)�Kv�|�H�`����}��Ǩ���l[@�j�D�¶�i� ��������&v!;G)�Ap�����O�̉O�s�pS
Fd@�D�����,�ţ\�M������J�����c[���둧w&Al�cף	�B">;�;A�|��5x��K����D�.�}�;�4Ђ�h��'���m�Y��!�\4;!�|�n򳖠G�S.�ݵY�j�e!�TF��kGgZ7T���|�pD�C�����0B1����Td~�歞K�x]u�ꨤ���.�gNT�]o�=��+��.���#	�)6��$AD�G�fO=Gį��'��l��盦\H5�]�7�7ް�L��:��j*ݠ[�bT��?�t:�`'��L���$�egh�~�&-�I��l
*Չ?��Ų�+�~k��]��qAc_B�!s�Èn�0�ۋ_s?�cK�7'?82Y�-xqW{-Otl�M��~`,��4^�m
S�3o�_�4N���(��b
#�[7�Q�=�ݗ\i8��_
2䰘��T�By.�T�R�(Z�ӗG7�N[�U��zq����s��]�WWy��^ ��uz� XGgB�-E.|�;-�� ��iq���I�#��#R�Х�0)���E�g$��_==Mo+Ղ���s�f�홄�d�Z��̶ccrj���"�0l�ȍ�C��C8��g*]ϲ�)�+��$��c����a.�{�U�	c0��8HH�+�v��-N���鬼o�E��%�L�{�Iew!��0f_��Rg�Ծ�m�!l+0�1�Y7�e��1]��u0��$[Ap���jj��ؽ~"OUWm2:`��V��N�������m���Zw��ܘԐ��=���G�ȁ����1z����	�[�3gD����*Ѐ�����I��JF�!c;�jW�oJ�����"�YS�W��J�,�^�#�B�������u�9��whBE�U��̯�j��(P��5�%p�#�#m����+!~*IG����}�j�8W���Jt1�1����⹚h62�Mj�EӱsU�8��p�ۣ;��1��W�CSF�4m��ڷ�-)�l���� ���n��R$J�1}���h�&љ�������O�f�#���Y�g
*��5��d�@ܴ^.�����)A��;v�6�=Y���{T_U����������x���X���\��7W�,�0;��Omp �)�$����x������oE������5q��Nح=��qxb�&7RƩ�V/A��s4�%(���aJv�N�)�1N�Y
ʪ��L���3��݋��e���l;w�2jh�/3Ԛ�K'��M�4�a�9u�D���R�+)SKc��AI�������)r��Y*E�]���@����R}/齩�����0����ϯy����c�J��t
;��Ϊ��z�9L®�- ����>�j4��UK=�Bsh�@=�,���'~�T���������צ�G�y��5����N�x����j�yҞ����"`BkR��!w��������R`v��ÏX�`�A4|���?����句�]%Zr~3٪2f=y���r/�W��h;�<���($|s�����c���}ǰ��[���x���Fo�fi�0.��K��
�(�+�1���.�Q�J(,�|�0�^�O�Yz�V� Q\0"-v��B��!�)�y0xXn c8K�z~��nm2��c[�u��������މ��5�P�7]����-����x�lՀ�[9�^hp��n��j8vx[6L���ҙ�G1� �i�;�#0�ò�"�,r'b�D�F?��B-��0�G�Q�m�]V�E���R2�HҠ4u�l�%���3U�X������HQ3mt(s�VA>�`�Ҝ��x����?Ww y��ܽ���R�����C%g������֯BQ[V��`謀S�F9��|�{��@K�f�-����\���hf]I��\�w��W^H�*�<�`�>M���\Ŭ�F�S<�Nj�K��K�]mvf�`���hu��.�Y�Uc��r�`�G��c�{F"ͱo����$�Zھqo�=E�ƪ�Fv4ڶ)�)��q��c�J�%����Y��O���T ��*K�3^.���F���]xt��':�3�t�cF��=�{��~	?�d�eXKf�wѐ�J�b]#�%v|�*��x����@uم��[�����V�$@G�ڱ�	���[0E�2%j�FyL��7KKr�AF[�������ڷ�k�\Y�����z	y���ƽ>طe�~/[�ґV�i�����✠�!�x�,F��^��^
(+θ�H�/���~� �o��zV��>�;��9��&X�m��5�}!	��I���m�q�9�?=ؿ�@�}z��PJF��ٔ�ĥ����3���nf#l�pL��8nzJ/���5�)hX���Ǡw���v-�����X<��o3,aB8H��hPb��@����}�H�S��٪���?h�S��43m��S����{&T'�n[��c��l,.�Ŭ�M?_�;�'�{��	�� �kJl���ɦD�{�A�����btʸ���.�1���"��.�H����cs�KI�
��/�������hH~.�#����,��p���;{�F>�ı6�KG[�D�8- �AQ9	+QOP-���7��@}t <h&D�BŞ�UӄD�I�<U��� ��#���R6�Gx�eJ� ��:�����]��b/����x`��,��|�0{8���eξ�Vjӑ��9=�;���v{��RE���)�<�ug�p�ǳ1DçF�u�9������<=�y��S6�2�<j�cH3�coYYF�-�+������4�WMr9�h
�?�i�㓋�� yc�ro~W9|Z�T��}F!�<�'�$O� zϵ�YO��t����e���a[���tЃH�T��r��͟A$:���"�"�Vf�B?��qR��/�o!�z=����d��j�+KI�(��
��6��D�o@�M��hl/$-6�QV0z�6�o>v�����fx&�b=fi�*U,��p�A<���,�I�0G��+fK)��?���I{�G�=�5�5��B�R�ܡU�8u4���^��x�s����"�	�H��Ԓ-(���*r��Ѻ�����Tla1aO��7666@��u�nh�ܿ�s2��0)�Gw���k GBv���q4��^��&h�2�k���o���[��׼fe�ꙕh� pQ�W H�FgT�dà`^�]3�:��q�\{�&�9ÌG]�|��6�Rg0���R�A�ع���/D�L��W�zy;���( ���q�k'='�g��:�\z�u�����de������c?���n�t��K�9��Z�q;I�&��;9�^t3	ٛ�Q���r��v��[>��ؖ1��w´%����>Q��1�K����O�_m�B�<�5����Nq��4�x����ƲJ�L��%!}��e[`2�8}��c�YF�d�@n�F�'z� r4*,-��%P,ٕƐ�{���ӽ-�K�oy���d@���Z�֩kj�t	(�86f��YOh�t�H�"��[Կk��h{��,5��~I�1%�Ԙ�5J�&m���)̜VƈF�y�>K���gE�X��|0��� ������F�mT��+�È�q�"�R�e[v�3.hLs�+��0�tW��F��
��u&�@�	���MI*}�aF6��,s��K�E�A�����Ӵ�k���Bf�֩!�s�&���t�S�.����\�[�r6�����]�~�N*���iP�	�V�r(ԻD�4�Qu� Gq[U$���ݫ���R�E�e�&㌰&1��f��w����%�(̖�&��yr�Q3e� ;i���,�[4 �C�����:A���9�&�ܐ>zBXU���2ǡ�8�>z�B�!���R��t��MNm�b��bl��K+0�?;o6I�����bT�y�$<�p򠂟1��e7�I� ̄�����_<wZ|����x�RF�Ĝ��,��Ւب �6s��ja�͐59�
��_]|�y(��G%D���!AM��
l#C+>���h�h���ۗ �3��*�rn�⏴�;o��k�}����Z-���Dv�2����B�L��e�l�Bs���R��b_qw�k���;���[���"&J�`|D&5v'�5nO�{Xǩ��	O���)h>��I�
����`���B�O � s3gѕ�}_�-����&`��׮�؃C�tp��K��:�N��LET�f��;�:�D��~�"/��J-��67���	Dx7���{@�7`A�t�@@Ɔt��Lx�����:��W|D博���vꑾ�q"l�+ɩ�7�U�,j�!gQ�A���6n��IC�-=௄�GM��{�y�[����&��G�=`��1�P˩�p;���\��-[t�!�boo-�?�����nt�pv���y��G����Ǩ7����Y~@x=
o=�׎q%ՁH)���61��ܐ�{�!_{������b7�j	��n�}����;y���ul?N=��fdQ%���K3��q��~nF=.�Q����U���
�C�rO�Fȸ񠿔2F{��-k�FY�P��� �K$�
(_Sz�y!ޟ�棭���[����)xR(�1ws4��>_'0N1��2�W�H�`��n�ݬ?�ҏ��:�Z����;./+!IZ�N��&�� DM��M��E7��gw������£�}�>����B��Ϯ~ �J��m�q8�u'͆[���i�G�7�נ�}�����A��iTp�b<��s� �	��-2��ow�J�KT����_�_��n=\4,k8x�i%�!�TىFH�>A2�J��2��������u`8J���=h���ɩ]�N��T�m&�ēkU��/��ؽuo�`j5���U��8�x���@�z}�9K�'�^0�0d�R�[�����:�9�Me�a��KT~g�MG����������D0T�'�ͅ���m�*;�C/���O�,bj�$��-�LQ�pN�5rp�@*]x�N�d�'���T��0�(�t�^l�P��Ц\MQVvz�_���hV���u$���3�7�o#����������Y��~� �x��?ʑ�w�$J�L��╘��Y���y���2�L��
�����\s?��i�$\�پ��u坏t�i�"�|���<��n�f�-`c���^~Rf�P�d����U�����L�õ1�-[HD����?��X�h��1J�����!�0�ѭ��ψ�����k��S��K����	�T/Q�����s�����w��KR��[�E��}�D2�y�қf��M�GZ�:Ƭ6N֌��"�F�dM��m���wA�#ל?v`�P�i�WWL2 ��'�Ŷ�'�e:H��8q�W>οF��l�鷀&��_ ��I�� �$���*��+ʱn�2fF�d��3�
?L�=�x��&wcAVחy��<�P���Q?9jJl���7�8W�$irߛ���'���!p��N�������^٨y��Tb�Ձ =;f���m�L�]f�E̢|���Y!��2h��Lq*O�Zn�U�;T��˲��-��N�5��Ѩ:����f�,ꑿ�1&}lYf������x�jx�����	!��7���E��_v�]u�bu�U����6R�To�W�����W�j���&�b0�F��՘	u%�M F:�U�9h)�xVz%M�R�&�w#N˥#k�����$�� ���@>M��`�+��B�M�U�ŭX�M�|!���?w�΋ԁZ���y� �����c���C��x
�>����Z��#EP�w�prnV�g��W�Ȟ�[�a
��hT�g΁yG�� ~*�+�(�B gK2zȑ@pl�B���X�������s��
b|�Xh�K*�	�RfY�D*�BnZZ��X��kN@��;ݪ�$����l��S�ý,	��#WB�K�]�1�9�2�d�̎���l�Μ觊(G=M��3�\*�]��}g<��}�o�}!%�ϟ(��S�ч��=NT�8L!��}D�,���ҲQKA���]0����y��'�v��C�p[&�p�ݚ.��W\=K�"���3�	H����u�2���$�-��<�6��qHփ�v~BO��r��Gkc�W��Y��#r,w�*@��i�!�sd$M<���$��l�}e!Gp437��6�&��]GZD����)G���gw\��!OG���{�M��4��u����<Uv�t�=�;[v���W)�b�)�����"���a�a�\���zZh�d@�F�Β	+J�<�a1�B�}��M~����6����CoH����V�_��%'hIF��ڼr��I��zV��d�"�|t>5{���e�	�u�{NB��+�:�Jl�0#�ȢW:���7N )�V}���gg1A����E>�l9�:l�\�k޸L���w��;S��f���`A� �����I� ̵��ڏG�R��B�d#k}�u�"�=
���r
x �4�I�����[�~5M~�c�	������q�s09��'x"�_�8]��gve�@�r_��F���`��q�\�7�� �[���;�\�A��{{x��ڏ���oӌ���n`����B��c�3����6�3���p8���a 
%��1���w��@C���b���Xӗ���Xo��������?�*���k