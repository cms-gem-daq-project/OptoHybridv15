XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u�=X:W��4��j�������
n���(��[�����D��_.�~�����I���<���9�sR����35ȴ��؂	D%�:�V����	�ITw0)�Y��� j/?L���6����ZbSA�'�`ύٵEJk�%!��IX|H'��$6r`Ao��@���C-�5����,���0�IK#�|���c��7���3p��P�OV�k�� �[��*�� IH�� ������(�@$~lRI,�۔*LTb禦��@�n'̃�H�1]%#�|z�ي��i�w��U�X�J-
k+$V�+�C(3[RA����Gn6#q*82s�ꊯ�jCx�#&�羳� ܋��V�e��i�Z�z˒?� �X��E"��Eyfb�^�	1�\cG/�-���.�zj����5��!�ކ�u�e�߈��9��������Qֲ�aڐ��]���3��׌"C Ͽ�������9��S��5u�̌�ل�����R+q9��[��s%*�7~We�K�ox"7�K�?x��E6�3����\S�OZӖ� htϨ��k���b C������mU�
H�m���H;jI_%����֍�
�\h	\NM�	X�+{�>;��B��kS��][�B��)ੇf�UϜ�ʹ۪�$�uH��l��@U�+k&�==�:O}z����(�9��I���1y�����a�	�z�eF���h�a_!��/eP��6q�c��bz<o�5�1&I��al�Vy���cXlxVHYEB    1577     5a0R��-�~��KC�$�cD>��(�5�-��Vy ���3�<&\����rb��|����l�|t@VW@8!�w�3��KJY%3�Зj�yl^��wKpv*�����g>�n盃X�^��3U��X���-���	��<ڡ�K�uD�:
�J��i� �����6P)',8d�b�F�����%;>��A3���S+ٵ��~G��.��80�66�Բbhׄ��X��s��Q�n�^�Q�� ¬|�:�4+a�{��;:t:�����E6�S��R��ma���y�X��&���o�s�m/�?Q`w�k!JqT )��Z2�s�K6�+���VAo��'uyDh�vCĪ�$CvS�ӹ�b�Źٓ��=%���#�Vh�}xƍ���ݬb��p�I>4���F�4��?������#����EFA+�
����81g�$��O0�͏P�9��r���k�<��k<z5��%��&G��c|�yd��W3��FppM�訵�n`���1Om����6&���&��)�j%�9����Ah��'C.��w
�)�6l0�8Ų�Y���8����]/"�x��ً������[&��X�6$�<Y63'�:��h��U|gP�G�)-j1Gq��h�w0:)� }i������z9mr#DK
`ְ)*���98�o�"G�*�}�绵hDUQ,��>�P��jذ�����R�`�d��#gvj`[��߰(h�j����C_���Y���Zj�k�����J0��G��N
I{����7�HO�V������1�j���1�v9{��o��8;[�6'���� �9����Y=�h\��f�-h
	�ϼ��m<sS���	��EUU�xmik�����$�+$�l,aP^ڬ���q�hq��1�E�;)�����S9עm���&�����A�5���,��|.����3뾠��U���lt��o�$����M=�P��������Q��=����x�	���/�ٿx]i�IL�U�#�S%N��8�/��'J�R��Ԣ�($X��6!��8A�G}��Q�:?C�>pX+�oy͚:�.#P/L矣#��$�d��ώ!L���������Im���}��|ծ#����'7���(n�|���M��5��1_�н�vj
�T#����u6
8��oq	6���e��@!�c�?�%}����J��Ot��Q�l�X6]Z�5۴9���Sz��&���X@8��X�۴I�l�5Ô$��E$N�f0GY�?�*@�Đ����	/y�Ŀ�_�݉9��v�	3W8C��>A�<\2�T��G����9��U��00���5w�	<d�=t��RY�t�k�bgOW�fx�ת��nypY=�DB�� �?A|��R��Q�F��n+��C��Zx�*C�,�i�(b2��%f��