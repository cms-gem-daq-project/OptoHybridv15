XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/���Z�[]9����h~���D#Gב�����0�F�Ic�W����ER���_�Z�=�����j:�M����u$�eiD���X��28��5!�i�T����-i'㗵Qد8�܇�P��_P�g/��! 0Q���������s������ϊV���א�����V�%S��-=ڷ���lz0��5���b�g�5�H��^����&��E
6HU-YJ뼵����@������5��Dwߘ����dOYٿ��/W 7�AВ/����Ƣ��j�S�\�X����=J� RTP������XB������w�̇��R��Ȧ9^-
�=W5���B���+b	�v���w�x4;�����k] ����\C�:w���N�($�2�����ެ�§r�-��թHM��߁�l�]uf��`�ͣo�� Q����6��$�n�;�^���T�p��>
h����T�;���;Ob�$¯�$;3�W�i�T_�!��ɵ�R|��/�;Ie�n�>��۶x�gZ�\�Ԃ�C��dǥ4�d�9j[�S��j�������)	�AD?��7�QW��/����7Rxt��!�t�,�h�d��@�n��؟F�($���R֎�v ��y��	��hyc�&D�������n�)����Ea��	��9HF�>4%Ȣ
����&opNr	P�x��.���)���ԄLͫs!����i`���j7i�	�w���W�?��Ƿ*���beYXlxVHYEB    60e7     cd0���S(�Yq��<~����)��j�:Shԕn��� � {qB8#U�>�,�x�h�t̳(�Ԃ�v^V�8�P��x�wn��!2�=�A �޵ӂ��5�������[&����Q<{/&Dn�ȩ��l]�_��XR��F����|8�TP�^'�i,[o��oL}��&!%*ц`�M+�A<O�^��|��|x�M��r֞��g�L]�î1��zқ���8��Q��;,7`��5��7s5�p��a� #�4'P�R��%�D�6�*��Ɇ۔�m����Q/�K�?�P��$!��J1�2'��"�'6C�`���2\��������l
F���� n�sB�15!��u�|�(�c��U$ۡb�"��+<���iE@�D��!V�/��{�|��/�����tIQڃY���o3n��	��U\T�0�L151�`SQ����9io_���o���Ê����]��*ݘ�۶�7��D�V��쳻�e�K����ݮe�$���ݒ�M�;"VJ	y8��J5�q�zw����O�B�p͏�}5����4`��*aJ�G�V<���d	���u��f*���Mb��:5�B�-ǚH����u3.�˃s�F�k�]ԭ|w۩�ŏ���V{*H/�����I������+v"#�cüV�&|E	.����󉪴'D8�׮5�O�**��t"
��+[�z`��NP%�Cƹ�i~��������YŴ���F1�[��t��W��V�UnJ�*��\�!��<�_��6O��F=�#2�᝟Ŷ�tZy����*	����&h��
�P#y�S����+�%����:��M���
�@_ ��"��S�ea�<�M�X��J�j��o׏	fXy1H��v����@�{��Ӄ�s�����}��
���8"x�(p
�:�_�a�x�d޽
�Cf	t]e����9��Q�*��/œ�F�����v�� Ю���$?3����8�_��$�;���N_gS�[+w���|̎=�Z=�S�ĕ�Y�큈�M��2��T1"[�����XF�� F�ჺ�#�����L=ָ�]�0�ᚹY�l��u�JS"��L3��s����� ��>G IlR7�����+6
 �H��/�󲱪s��`��������Ѫ%��Эe5¤����n|\�/��Ҷ�L)��S��={�dp��=dli=D��]&m��f�T�z!lϪo=�������{j�h~�*�>f��b�z��O�p/S��p[��;j�⠈��48,�^K�~���rڥt3]��AF��؝LJ�.>����o�'���<Nֻ�8�VCh�~��+]~�<�On�:6,'$@��fLi����I3tqnb�
��6���nɿ�:��E��0� �[��۠@K0����Uϧc��j"�خ%�:����%���Fz ���N\nW�
��Lc��)Jv���,@0��q;1��V�>��ͯ�0&�4�fu��$��3�xj�7f���u��!�$���RF�_3s�]�������h}}KFx�S����ކb��F�k3�ԮϠ�c�e�A��0@��۽���&5�9��=��Lrv��w�habkS.�4��f7�Q"XK2H�ϐ�]Nb��<�WQ�]�\[O�sݍ�}�O��D=+=��2cÛZ�GY�1OY���z/¹?���y6�ҝ��s+_��x�N�J�7�ԏh��9��?Lҷ�]�%�RG�����/�^�N���Y5��cK6;:h�!_��e�!o��������\�{}?�M5��.*ʊ\KJ3`�?E����~v�X.�
��Dn�6@�~$�rn|�A�`W�87�Ti'^@6���l]C����wc]���D�5�h+��!#}��ﭣW��.��s��/H�.�1C����7L��N:Ou<R9x��D��sx�`d<k�&/:������]�C���Da\9���1��ms���gG���{���^�m�Y`�_|��[h�-ή�O��@�Rq�� x��t<��S��A>�,���ճ|������������U�8+,,؆�$�C�B_��9Z�!��]G;��H��k�[�����8��à������2��A�}ƕ�c��4�vKH�r�I��ޟե�9��P�ݏ�!Wb9;nN4��\�$���[�p �C�{(Z�U�Á�%HU��n��	[(j*�вNU�����Q؃@̇���v_@���`����7�h\�')�������ώA�}��3u/1��m_dk�A��O�ٱ���+ݮ��f�^b[)���s�_���?#���>�1d�е ~�ʠ45�1�͍����э�	�Y���l(J�k95�0�x�Q�?S\A
zU����Tiۮ��厹��;M�x���������"l�;��[�[4�!�Φ#�2�X�!�W��q�#���Q�v�E����Z#�/�m6�����<b����iz��� +��5�jU�0��6�	�~h��8��50ak�"�:�1b륾s�����
�r֒ESL�w���(��&��;u�{����)	�8�n��	쥥ec�%I���KdyO��P���Ѓt�ޭRX�C�6�\|.��0F�v��QEJ�+~zp��8�L>d�+�l�i�;6� ��u�!���_�b�@�U�7"O!�Ua�`��SA�Ʌ�pDt�-��H`��__bu�*n�M)|���T	OAY�j�7��;��TUz�H9V�dz],`�լ���f�����'q�Z=��C�+�������뤹XV���u�u@b�,+�K滮�����Cm\�-r��O��v���8����!���E�.���1�|ٺ{ �Q����_�%�>�#��o�6�9�X'����$�О0�7�m"�{@�<�AUh��dCS.������S��0�P�}����۠��GO�Ð��2��g+��=�X�Zl�������H��I�%h)`����Y�6���4��� E]C"(�f���6��|F�BMr��%�܆��W	Dq`w)U�䩒�j���R�ew�/���D�Ͼ��Xt�I�<�E^0��Qj��hb�#׀�-n��Cl-�)���g��!ߝ!�'q���w���HY�Tr����n�d�X�
�(l:@(S��n˓5�	}؋�[1d����Ie���t|l���h,4f﫽�t��2]ֲ{�b��#~r�NN+z�V���ظtw�f>?