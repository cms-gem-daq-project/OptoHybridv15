XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G�;�aU��9{��l�?�<��TmC�Z�cd�3z���g2@
Z��:d��6��.�vTX�[`�v�'���:&=	Ӄq#�E�q�5�H%�
������h}���H1�{D;df�����;��L�7�)�zd��%$;vo�&L��늴��?��$�	FC���U��Nz�=�SE�R'�V&₧�B����zS�{d�0m�M�����z��x����	,�^oA�J@v�6o�h�i �x�XrH��S�����D8F�#�˜�������M��Jc�xFD��>6;4��!��������~�Y?��˱))���#���@���{(�J�d5�C��+���Epu��a�FW���o���q'�����v�W4I�F�;4�ULnF��������a��%�����50�򾇫����"7���tH��k������)?Rzx�x��(��.��� ,!ʞGK��ӱ��v�S�%
��Ð:N��R�:��OU>+0z�Z�Τ�o�QjH���l��F5%t��KK�p]L�@�
X:yİ�i�.���ο��Hy���~Sk��,c�8.��O�t�H��.UQ'- d˧���&�."�v��l�m�u��Dg�1BĺO�mK]̄¯��R��E��U@��y�M<�ϰ��G"G
0e���C�,٤O�0E�oP��|(+���_�������e]I���fЎ,"V;@����I!r��
�O�[�h�?}�|�u�z��jXlxVHYEB    cc3b    16b0�+C)h��Z�Vym�L�a�dE뜎�-%(4ZK�a6�=/C[�ҹo8]�ܴEV�[XVi!���Bs���W����ѧ�c"��j��!#�θAm�� ��h��O�X~sbl�i;x��9�g��w+v��I��F��}���;�A�&��bЩ;Y�֤5��+u�)�l��s�}�c��,�Ud�u�c�O��� �\�jb)�o/"fj=�B��B��w�c.ay��M��4�<x0Gh��`'aװǁ{ֶ0��4f�O^{-�i^S_,ϼ�l&Iq�Kƣ��S��!%gi�&?x)�כ�>�Uq�Q��s;�Ǵ�E;F� H�p��o�e��t!k)�*�Ogi)��|W_�W���Q1�Wyt�)�Ѥ�Ѻ�)Ux:u=�nE3gi�ܚ7r:^���V^#Y0&����(0v*�`Kyc�$��%��rR�;�ȿп)'D �m���a07m40�ޟu�۞�{���Ct*#�a$���u�����!���#c�gțB]���1�c��-Ny�ʊ@�#2*��vE���#�<ˀ䒄��FY�z&iq��R �4iy�jO��'�=W����E�W?�I���"3N~�j<���7YtOA_|�G��-o�<Y�����i�z�sb+�8�% S����n�����dec�'w�h��Qf�^v�s}�����2�=��'�&��3�ڬ�L�!wN�h��x�Z�Nm%�1�y�O�Ӻ�S�����76�X�qG�O�i���GZ$6M/��9��B_������aT�ҍOI/-�Ϯ)�C�c֔(j �4�V�ګ]���v:6���k����~�f�6�G�Ry�)�X���5�CL��iҲ��C�_�	0t>��54ȡD�s�t��c��(�wFs��j��i����7x��S@z�A����������i��K�+'�W�ت�!ΝI����c	���Ma��3����t���Lԑ�)�
|g��1 ľ��ܯ�\��d��J$��ĳ�T��?�W�^U�p$�`�N�_1o�i+uF����_cL��z9dh�&Z>/Hv�([���;�䌚��z�+��˘1�������2����_�;����&����Ax����s,�ORks��yy��챿67�\��޽L21s{�6���s�o�.S%�ʭ��F}��$A�C��'2��a���o$�C�Q�	�Q��7ψf��[L��	�i����o��_0��RI~�;�C�V�]�~���S9��@�`��V)�v�7�0>i� ��#�w~�q��ÈmTw�����s�i�'3֬�D�C��2|�^���c}�5��qd�2wj�<�{�	�wnT�U��n~�N�����2��V�cGi�F9� �Z'e0���~����m�|���}���D�b��u.g-)	��Cg�/y�=�S���Ě�	"̶d9�e4�"*5�|/�nF�SY�8��`��*�S��"8���0�6mG����l��(�O#�F6��+���M�\v}i��4��3[P�U%��R#&ժ��!�����3O�ǫ1����_�-�`��Ϩ�i���`6�ޱj��y���B�C�x7Ѵ��z���L�>+U�׼S׳f��_�:��;�^��o�@�@@�S
�>���Ϛ.2v��m<V�{�Sj�H�Zsh9K�<)P;�.ӵ�b	���YE{��h 01��C�����ZT����ozoߖV����*�a�_������1�U�L�Zw���lB^�$����0nO�<�Y�:y���g,⊸	�X���t]����G`owR��j1�Ki��?����l��ղ�!]��Vh�Y%;�����D��+�Y�����!�t$I�d�0�T�6a'�6�hV��R��}e.�I�Ƶn�yG�`;���B���/F� a�����O�ύ� #c4�������p��j�����
�I�$$�^�}2@��7�ܣ
D>Z�:�r�;�ș��(ho��5h����X���6T`�avm>��GV8 �R"��������t�7{����L�ճ쫴�}?�����P��C	*���y�^�������8j�^��̋���ۄ;����2��4� Z�j��J7zNO����,�e�<D��`iS�U�\�k�4���l-P%�eg�嶗��{Ж/��O`����>��D�b��w��+�Ͳ��3�BU%����֮�����,����b��<b�B��/�����o����6�Nr���_]�g��>��N��w��!>9M�p�ho��':���~y��:+f�lyS�	��^	��2vv��Y[z�q ��?�F���1o���.N�����e��|�^�j���t�f��Z��2% �¿r׬i{�u�3��6RTŗ303�*K^���:w�ĎhiS�9��!�w��*HOҌh�Iv̞�,�Qc�Ofޚ℟�
��뉍�T��Z�J��㇀��<U����ѕ���}���� �%��H�� ��,H�m������2����)e�4S����UY5��/��vsfW�TPgǍ�W�tn����Q�|��欗�4.�ier}7�O����P=���t+��-�#���1��|�h��9ط���T��;��Y��"�&4�5��@�!������Ap����"$�Q�9��V�Ğ�M*vr��4���較q�[:�1���@����]������~�o�rzY"���t�>�����������:G��g���>A����.�O�c�i9�D*�-S��/%JM�O;�"�T.������q��L�.^�C���`�b�3�W=�u��
]�cg&k������������rQ��hT%,و7g���}ݠ�a$���-� �����=9�P��r��F ���]L6�7��vǮ<P�)R�w�A�4�5�\��SE�r�,d��ca����kV�����H���5S��r�4,�G^#�~Y��'�e#������y�I7A9'@����2wJ�⮂�Lu�C#�I^�ʊ�vs4���<������H��0�8�`#�F�,L�Z)`���G��Z���m4��E ��U
�j	�ok{���N�`d���آ�Q�!��0qB��Q�hB��\O��&��2�V�a������<:��>20�A�(���̛|t7�ɵ��u�5q���Ⱥ\jK⇧g���-����P�M`�<kFO�����)4�}�TT���#_t�3�i�K����,:��1�&�t��.h���Ke���קQ��>G+4�8͕@�A�E�b�%r����*4�|��7���h2���Oth��m��uH�D2�������D&���QJJj��J�!4 VOo�l�!ʂ�G*��.AL|<qVw+�E�?���6���9"�J�w�e#���)Tc>���UQ�?�����p� �j�1&o4�ccWk���>���ZN�=p7�4�0��� |+ZR�kY+��%��g��@���:��s�N~1�A�e)���rR[��Jo6ߩ������F#]�1ǒ'�Js�Y���겎 CiT2&���ǎ�+�qN���؈J�_rb��3���D�#ׅha���v�Ԁ��C�*h�-��,wqY䡍�P_9�S�>���{�V��x�:�W�����:�����Ժ]�97���8����E�
�Q�IQ҅�}\y�%��Q���,<�z06xf#oY�C��X�;čb�-(ˎD���>^��2!3�{�tın��b�kn+�0���yXx9�Z9�P���z���y��e����N��D������U5.�ioA(�Nz4���(�u��-��[��a��-�F+�Re�� ����.��z���l�����CZ.t'��K��و�Q�1lVF�ڻ�a�]]��`G/%܇��� t**U�C�Ue\ ��z�ᣃ k�Q:�)�A�}�>�S�H�9]���Hoi0�\;0�uQK�aN�ܒ��e_k�iH�G湮��W�� t!ؾ�W�ī��o���ܲ!`	�~��jr+�|��E��TD��6A0���ώ��x��cã��u�`z�n"s�#�߃ֳd�E�pq߇�.��؏`UM	�g(�vP��S��Hg.xd�;�P�]�,J5|�A���# p	��ݴ�C����VO�c��tJ����'�07]li<J/��##Y� n�z�7��_y�Ǎ�k��\����x��M�Ewֆy�n����0|٪ES�ꭦ�$��-�>�]�7��"�i>�ϛ�R��T��0��&R�n� cʉ��ٰ������m$��e
aǵ��S�QL��wo�L�*J��_����$0V����K;ǋ�YX"Āri���ۓ��9.��U�*���P�c�4����D�nI4��x�k3�x��	�qY�ټ*���L���Z�b��Z�Ndwp����X�6�*$����1�忳�X��*E�M\��=�ޮ�"�<�!/ؾ������Â���w�k<j{�u�nH�o�$�Ӱ��^�=�k��7>�l
s���3&ԩ$��c�@�';-n��w�T6����=]��m�b��
�o�s��z�W�u�w������{0��4M���̉�yq����6z�1��m(�<� w?L?[��J���ڄ:c��Mǳ�%�B��+�^De���~+�I�Lr ��1H.>�zU�)�^�p�����_��J��#��1�{z�(�Z�,���&�rȨ2>��6�����Ǚ����I��Ɩ�H���ȣh��#�xo��b�{R�����m��J���R��wG����XkVPE����� _C�L�� x�;��{���)���d�A���}��_�Ef�e,7G�ǲ�a���}��$��Ƽ�l	C���p�b��=���f�� �<@_%�xJ�>��y����n$�y@�zS���FLɯړ����]��J��x_˦w��Q&�dk	����Z���֢Ғ9�����.F���џ�HBɔ���vn��lP!t�Q��^GPlӷ�1@ОZ�f|�b.I�k�a�M�(�]UiE������Xtô�H5
��7�n�4��o&��U,�
�����j��(io���ȣ*���U�O��|��t�4��rWpg��Uoa�T��kS����L��G\�4˔827��nV��?y�GT'��)�Տ�˜�E��}t� �� T�d���6z"2{��r4�+���J����C�v�c�8�,�%�1��� ��w=�#�Ѯ3 �G�&ҟ$m���Lg����A+'�q�z�mؐ�W$H�V��ղ@%t���sO1��Ïi%��V|T3��)~����O���[��Ƃ�R�4ݱ�`��a���b��Q	������#�u��w��I���Hl�S&d������[&�\��� ��<7��)u�1�5��D�"*�~�@:�/�o�
���x�:/B�5��e����+�k�駱����A�j"��a3O������������;T:�]�n�O	��������d_F��9A7��25܋�����q���N�Lۻ|�T�,��K?�O�ùg�+�z�|�K��u"�'O�j6VU�8ʵ��?U'���w�	��Y8'�8��t�1�k@ؼzS<S����Z6��#V։��)9���*�2� ��2C����N���D�d���T���=���'�ن�b��z߾���ڽ����wb?�b��E'Âd%�u��z�֔���$�~�X��h�$`<���п��d� &�Cf�ίt�'|�H.���