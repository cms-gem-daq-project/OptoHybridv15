XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����V��bs�L*V�%����������8��ʨ��M�X�[)�5�6�W�{��U�{jV}#f�U�����q�p���)Bu�/X)������6�^1m��:��2�g��������'�R^�)򿮿i{N�A$�q���_�s���XR��>2�%��×�zC�X���)�KNC���U���)Ŋ���Gm6�n=K�������W�N<�C�O'p�	z[���bo�1��w��M�:s�����+�M>�[c	�U������'X�S�$��8�e$���S|���	¼����I�(���@�����������P������d���m�2���@� &HW}�H�(	BEk�x��^%SS�[S�*���NÈ�F�|�N0sR�,ģ��)��	B�t�SXRZ
E��G81�D8�B�����+Y�:��*:��!ű��O��@)��_V��l���WdR-��I�v���E_	p�[�{���Q���'���O�^��&���f�������z���U��zO��!�__�9��a�R[$�X�X����?򨲴i�5��O`�S<K�� ڴ(Zx)����7�J?W���
R�3�*dmB�t�Ro��kN�j��1��"�=�`Nn24�I
���V�q3�Ō�]��?Vz��2a�X�G�x���+�YֈK�	P�Խϰ>:��p�����8�����5�~0<�ttĤ;�!یBq�~uz��U����_�W�]�4-#�l�
�<�����H\�i�0���XlxVHYEB    27ed     8d0!�6���MB|�F85�yI�D�n~��MŲ�!�����PdWC�!R��&�6MK ��*~E��V=�{3��_RTD�R���W�S٠�S�x�Mv��m	��AeGZ�5'�o���?czy���6��:�d�`>3�d��Ͷ�"G�oxhgʆ����+N�,�s�9 >&�zd&��yv�Q���Y�7��2j7e<�u�{ E�Y[�.r�!��=��v�t��u%@M��\TL�N�[r�C{|�"��Y���p^;��"e�I�r��<�ͣ��t;O� E��?�r�S�A�Rcy��|v�:�6w�8��X�_G=�On�pM�d�悹��'�uub)��O��>H���a��.m��I]0�3tY��-H��P�>J�+���U�K&:hqt��
M�)��/�k6/BC�2J����&�'�@�v�k���H(\[�uHZ�y���ڕP�����w�/�\q �����|���p�\�ڦKc�F��R��������P�� ��A<R��˂7��I�lE��s�K�e| ")���e�Y0��"ȥ�/Y����MRa9�n� 8��h0����,	��L���ɻ0���O�H ��ۉof^����WE�\)r�l}m^��QJN��]�oT��}ة�]��w7�a��T�T�#C�$m�)��k �}:6� 	��aM6+MVߢ����!�k��82dH��K�1Lk^6\j%���I����䱆��F7ɍ�ցJ�|_����8���p�{~L�Sq2��W���&���wR���f�F��î-Ԯ�����k�|�Wc�Mƈ���Р,-
G}�SK,�B%���ô��VaLa%`�M�Q���x��T�"A&�!�Km
!�L�=�l����Ԛ�g&5Q�v� ܭ%��)n�0e���*�jƮOxt�&j���(��sRn�6&O��TC���4\�}fWa{��o�4j+��^�`m'�(j�C���XrL�� ?=Hz��w��w����k����Tsξi����!����<[�� S��&R6�����������٩�k�}�i�
,��d5(��%q+��=p������k*�t�#�zϱo��q#8NDd�I$<a�V�O���K�W�a0�<1�|M���C�zl��%W�Ӧe�ьPd�雟a��mlP|4�it3$�B�� K3'y�ի�鷲~���_I��u�@.4H_'Ha���%~F�cf��H6��A��,�<+���uoO��?��j�Uʢ$xn1��Z�]�R���q7>���y+d3[M�`�_�9ۉ��m�qA��I�{�Ȥ�6�n�J�VG�WP��n�G�ح-v��8��Zy|]�f�T���?�*�$�*^��{�jb���ؔp.C�	��J����j�w�����ا�gb�<{�'��c�8�r�_��:�od�7��m-}b�rӞ7D��.��hy�A@,��7���}_P��Qo���z�T�gt�3*�Vo�D�aj��3t�
d��-�a<�[P���.4���g�]�&V�����}������*U����bx�����&��]+��`�_�Z8��֌�oU�f�&w�O�&)�+Z����8+;�B�:W)���ji�62G!����b՚;�2�{�Ŗ�hd���YX�!%�xG ������h����W��X���
���+�t"M��n��o�kJ�k8j�Wu'��cMǧ�"����-�Hg.>R	I�4�'�/C�AY��;���'2��A���!�T)
N�����y����{d��_�鈢M��U\z2�N���A6�8�h�`�*�N����zD����s�։�WC)
�;0���4Ll��"1��J�b�VE�L�N�%wo¬�~�#�b�7���訓��A-���DH(�7q�-�F�j��'�Yb)'�l��m�,���%�����?��� F�(�զ��\�i����`(� J��+��H0�C\�*����^��N�u��oWn2����.�>.�^,�Ri�c9aK��$%�sEQR��±���L�=���@������B����(b/�_N����?��ܟ�QטDe��ujA���v��#Yu'�TF�169�-�����㝱J��'����n\�X�;#���s�;8Do�"��wK��ɹ7�8"�h�6� ��"��\�=ɥd 5U)���Ɍ����,b���