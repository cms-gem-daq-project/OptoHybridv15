XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-�X���Ŝ|��~8�cQ{?�	ڰs>؝�	6>9xɖ!@'�BZ��V Dg��U� �}���n�n�a��~�����T���J�p�Œ��Q��q�/4L�RI�{����Lpn�4�Ե0v�LI�v�U�{��S!)��PafcK�4d|�Z?n�Bk�`�e���c(0	���M���J+�d\* *�`�v$g�!�/O���({�s)Obf����ݻ=C��NE�t���3I �u����� ��W�P�A}�[v+�l0�w1'�g������X��&A9���AO3�Mӕ�j�W�B�{��Wɔ.n4(��h�_��I�ڊ6q��܀�t�,v� �$�GYو�V�}��n���)Y�jF��m%>�R�\����y�mY�c5HQ-�x����t��w�?(���K������c?�y�[N��֕���>�P,�+��]���X)��֜�"&#�$�<���Lf�0�HƐISH��)1�=�@ I�y0Ov���A8��ʙσEэ#�ҕk��J+��2�6��[�6ݏ�� �?���1&ABUB��z�{.
��4-ր����4h���a� ̾.��5��jh�t��F�Z�6�H^���U�ž;���͙8P��ʌ�����Y��N:�%u��ʁՀQ����t��|�Ʊx��C�Ɖs���	��'��H*8/�̒Xq�y���V]��n�T�c	�D�[dl#�Ͳ��Wl��	��
*U��Z��Z5^M	l1W' �X�.����A(�3���oXlxVHYEB    41c2     c40싅�2S	Y���!�+x�xp�UBlI��f�Ȑ��[��7SNv@�9���
Dt7�ǟ���Q5����CF�(i_2�X���c��N)Ҵ�̈́�	�w��bp��1fvG�'HU��r�|�j�4������d��
�C��'"��˱��ɏ=��}L����:����mlv�%�p"�9@��I�/�%(�h��iFS���E���(~�_~1�j��e��xqMl�\X#Wj�/��Db_�ʡ�y����� �]�����]gb�.�M\�hP&��կ�$�B�U�=|3�hk�RGf>��uDK�������~Ć_ƠO�3��W��Ѱ�0C1�o?�^���o�SͶ�5�ș�:"�,q9�BѾHPZ��Sa�%EH���t�{�;��sǺ����s�:w���������А��SQ���:�)��	ݒ���3�,r�&U�� xUT��v#����t����P��#�G��� �~	��K���6	��ڒ�����N�"���D�iKL��=)�%o�Ç�58��wR�[IB�C/x��l ��"_+Y ��ډ�;��ȭ֪I�vW���R�LWUg��cg���Q	*T/��e�X��)�w�������ff˅���FZ����G�C�Z����y��d�&�33��'s�Y��C� 4m*��ھ�o�"UH/~ߩ4���n������Dju��Pc�sT�1���
i1�X4�7V_�諩�b&X&���K�c�[�[6y�-�kLjIڃ�o&Ѕ��/�f���P�橪�=�"8��+�fL�@��`��W���6Ă�(Le:y�P7&����6r@�WFT4 ���d4Lb K�Eϥk�{*�9�h#f�[���<����R9�$eYRjf~�������; �ً��ʒ%��e�< ��#��th��[��J�寭X�����줰��v]�I/O6��'��b�;ko�{5��s����t���|i�������*ec}�����T�R�@S�g��y�Tz�R���V������a/_kJ�ޡ(yY�'Z�&r�J�+Z������`�y'u�i7�j଎��)�pV~���1��ږ�O��/����}�PT�N���&�ud��~��4�)#�;̽���+V�fC��v՘�-<yۏ��=h1b���Qf�!g��]�P�?��)�����$<�T.�9F�$��3��z� 7����_����.���a�\��B�}��iEb�fB��m����i�����${��x�z�`�=�L��'����ðMZ%_.�	1��K@���ɸt(��~���j�ٺ-����B��pX�#&o/�V�\�Db�e�V�_�p"� .����+��
�[�A^��f�����ř,e���Ma�ꦷ˒�zQ���G�%��nk펨� ����6췅����x����`�tMgc��ӗ��}�2���)XW��F�l/��ۂzy`���F�x�CwK��U>s��NN�k�]$E��_�y�M�=T�	;0F��(��+����h���쬰}������X�v��w�h2�H�-�U�M�_�rda�y�m�|����7�o�;0�8�v�P-�={#�F8Ӆ�I�Jx�j�F��u��:�]�r˽�Ѻ5� �}�&'nR|6�-
>���A��C<��Wt;%�h��Ej(�m�O"�s���)�n/����{r��k�����%g8s˱�����NsP�@�W����<�i���{3 W����k�����W#�g4����Q�h��)�%}��͖��s�����K�[��������gΠ��%U�r�)��nh��Sn��掌kS1�� �#�k�x#��C3D�$o
`��6c�����c���G!�!�)=	OD��+��x�����E�z�A�)%BN0�4�ae�U��*O��Ggن��D��Q�.�io����iK�6��j�Lrn�"�m�����rkqR�����Y�ŝ"�=�M���:��)�����`	ݢ���q"�s({(m�X��VS�|�0�9�Ʒ�c���-,��\����(��@��>ó)]:gV�;�5���&��/�}h�ߪ�7���Y��ByVl%�`���uf\*q�jKL��%SH����8�����k"���o�B*�� ���nU�W^k��YN�8[�\[��NiC������˥��Jgmn�t�9ʆ=,����`�#������T���'�4���c�=�C1�,x#�^#ȡ����_Y=G{{�������u���j�?�*"Ep�kM����H-l*ք�=c|�1=y=�w�	u����ƣ�<�
�}��fWc�(g��`���=D��°��Z�q�:$R{g��s��Nr3�@�K�1���L��6~����0p�)Uz���^�4�q��G�������W�g�R�b!)�����+QO���|���Y����P��&:�R���H�d�lql�p����~�w��.��6q��|M�:�]?xp����x�ۚ���ķ�n��U<�:O�\���(]���y��`�a��I�;qDf��/͏tcwD�u�%���]m<_t�*%�be�$r �t��*�K��=C�rl����I!k8�4�pʀ#���p���\�EM0�7Y�;���V�w�Z��f��GN(%$�Z��S6.���X�&p�v��D�/n�����#�-ä����?��ֺ���*��`2_���^�-�4I�u��"�G�ʸNkd/C�>O��s�?�D�8
8I"��N�U��¥*�BUႏ���	E�"l��U����,L��'���G%�&3U'7�Hj��dfĲTf�pK�T�Y��Oaۭ >�ܞN�v��+�D-��m�i#d�eԽ��W�jә���K
�.Hd���j���Qi�WTC�lp�J�K9%iZ�1t�h2~	FY��*^%3kB<�����h:�J��}@����Dn��g�L���f��Oܛ��:�4�%u���nI��+��;Δ%ԉ��-l͗�Z"�1�կ(F�C�{�XHQO!��T$��V�o0�)�E,�r.�Lw6\(�V���)��Қ�j�I�c���D��|ѓzeT����j�����=�