XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���l��?�E�����1cZo"��Dl�򬒲�ħ�}b���T~Sc�MU�P3B�Tm�M�yDG]_|X"c�	b�0�>�cS�Q^孎R�R�֨����.��� �3�H8b�4�0-n���z�>������';n,�:|���;����p��ҦI�u��N/*�3�����gW�./�)N�����Z�%��̲4x�j�N���%��]��'�"��n�����%��?Ά�Q��Ye��/�ѯ����" ���Y#��r�����P���7��}9wб��=��3�S5^J�.Xy�*���gk�=��0��5��R@�t~(��fwZ�?��r���ɉ*M�c,ķ	���M!�?O�W{Y�X����{�u������o�g!x���Ů��a( +6b����3�2S"�Y�?ہ�����38!�;<w��t͐�]�XP%{&��	_?�:@���PՈ�;'��YB�
_����?���a���y���[7�ݎ����v���D���܃����G&q�geDw�U���I��.HC`
�uB�_���Yef$���� ��9�`�YW�>����2����{����!6މ���"ϡ��?ϋ��-~Ú�v��"�(�c�!Er�JϮ��fV	�*��!���T�n��&�1gJa���~��N��yV"�N�y0�rK{B~�J����e<U50c&����W�4���X�*m9㘤�g�>߅�3�R�F�v��=�6uY��Oɯ��sXlxVHYEB    fa00    1960��~�4r��87�+�y&W�N0(�V��/����������B#�t��)Y��Л6�s�밭���Фi���Ȍ����M®}4��´�!���Q�������W�(�}/y�ˉ�!��:ai�^�]:���ϗ4g��|�� Q
�W��?�$ug-��^68������k�̡�R2��9^�qˁ̐�
��.e�&� �TQ�"�F�?��vZ7���05����w<;�5�\+0o��d�̄����e�w?��y�@�)/��z���E��Il�Ypރ@��K��ΖKa��~b߲?tV%�*���������`x2�T2{��*H�9V/@�$F��`Sa����э ���l~�,��(U�a�X�k��5K���r��|�j�p�@ f�2�h`�U�]JhU���Q��nR��7q�uJ+B�%^�>�Ξz�ϼ�wU}�6�,p��<���`dM:Ex�vı�"I��ef�{��mM��X!�A�[,d\�2*�$��C �+��~�tHVy^�3lW~4�*In��}E�,��F�����hQ(>t�+,)2x�j�w�m>"��u
�h�#����w��FZ$��%&�2f���R��jb�5?g��&�L�w`2��4�I+EKl��ę��K�J��OP���qr�
Q�&�Rp Nkf�KbX����Y0!rS���0���F�@��4�B�ӖPW�x@�F$�żl��?�J�d������a��x�y_$r�qq�����t�rY�	<���;����fI׋��Wd}GS�8K�9I8�ri�N���������`v�k^f�c���_\6��t� .9��gkP�i��oo��G3�!JlCD�Dמ�!P�q�N�������vi��/v{����d����8�o1��A���?�I6Y�[m��҃"�MB� �����G�����o�+�V�<�$5�*uf��"�\m8���J�6�I2TO�xg�2SYx�}�i��㓸��6W�_�@r�РrU���-"�������26'?�������q�>���YǂΣnֵ��gh�x�?#͙�7ݪ�;���q{�%�@@���?f֪����ov�|rgo��e)u��S�\
"�.�?�esb�}-�L��TҨ>\H���)�ܛ9R�T��`~�6�T����O�=��U�inJތ�nf������}29�J��7Y��t!V3co~��B�|�0_'�^��	z����i���[Sob	�P��n�E-�x�V�ӡ�4�4��y�8f�]�����ΑL����T��7&�-\��u�N�3N�&)�����o���KH��L���#� ��$��E�n~�5qA��#�=-ک���#!�����aN��>ߒaY"��1�7�C�ׅ<���E:�y-��?�qz��5���`~"��im�*e-�XDV�3���`�*�ʘ�.�ݍ�2>��6qT �g�q-�u;qDaGg
����>����9_:������<Cп��\Yy�T��/�ZSdjw�@]aׅSW�=@���{��K��X�K|�^˙�9�G���}�1���a�g�-|;�I�\H&�	[_���g�N�d&�r/�� P ��!ҭ@7ׅB��+�S'�����Ʌ�:4�c�U�N�a�&�
�o�3���ik\�1�,�_�b��)�6�x�j���g�ng��q ��~��gڶ�y��{��&��ǏV�Y���:�bţ?���&}TCC���TI�˄����F�+�.,<���Wn>X�[������ -����3����B?6�M��*�gT�7�I��o���Z��<�Xgoo� n��	���n�R	fa1U��f|&H���s;}�W����D& 
��&���*;aQ�&Iy�!��n�1G��@-�3�811腡D`�Ǩ�R?j�8��?�(v!S�NG�2WS���P��\���V�j�v�x s�T�rp���t��ǆN��P�wDÉ2)Z}����L�j�i��+L����{�k�m�3����ިYZ����i_�k�P�;-'2�t0��7��^=Dݐ�����Ȩ+�D���nḉw�
3/٦1|Z�R�$��1�s-h`�.������C��qG�D
��bb�6���w��Ӂ��'++�d�:��>�@�p������ꕿ@^�or�W��$Rzx=�)�9��6�!�D��or�0�jP.����$����Q�(�$7�RQ��|:Lc���ƥ�4�y.X��t�>�M��@��w4�ʸT�!92y]P��_x����QrJm�RP.�� ]dٱeڕ������1��)�p�D����bz���܎�v�h72��ô0o1��>��g���x�Q�~��S �����EO�,����%c�X�ƴ8�퉲�ٖ?�r>Cܽ�u^�c��jS���#j�����h�$��.g�_8�`{6+i��P������gdN�R�Wy�u?%���WѲ�[ډҟ5�D"�p�b��[V�<>�,Q���+���LDX)n�(�׊����7h�iR),3��R�܃��Z!'F�J5�Ca�B�g�)�����4H���RAj��^1Rq�#��9ܞ�69�2��8��:y��wݐt�;����$Η�T�em����l)&��%��2���;��f<^jU,x�|b�>�K��^m�m��72#�&
�K� ��J%vom�{�u�7��.�q)l��ۖ���������F�h��U���ҳk ɧV��������`��q3�31c*�J@�_>Q�E����R"'p��W$�Ng��z���
�T3pv�[���ƒL7� �|'��om����֊���c�v42�E�S��f�@�t�]�3wIE��~a@�r�/`|s�A}P6��;e�PSh'�,Ρ�Lt��6�/S@��lh���� �_W��X��߂)��]���s���\;[��(�{�i_�����%C*"t	V���7َ���o�7�u���L�2��e@��*���^�F�Y�2\�R�� b�(`��:�K|<�X�o��;GF0�㤂2�Pr��l+{���ݑ+�R�C����gd��e?d� ���aG�s����-��MS��aa���e�pWZq})��=��%�2B�H�ӹ5/��1�M'C�/�����V'�d��;�/_�+&Y&Ч��e�D5�X�D`��ʱ��pHb�\rH���P�=�^���=RJ�\�1>t� K���W�����|VD��5�G���U7ڒ�֍P�yY��F�W����m;s*i��d��L�V���z�ґ��A�c(��=S��1�F��:l�6Cd�#4��g�w�Hl�F�	�^le�W�/�yB���2H[�_��X�#Zh�E�r )�H��_�q�|�s5�T �����K�m=Ja�:n� ְ3-�#��A�F\��K
�-����}		�ʹ���H!��|�-!��� 
1� �:p<��>��w��4��M�.�s�v�W##�m��hHF���p3C��R��������v���S֟`�zN�ab�=` |�B!�$q�ACF�"�#���Ri���T�nD���-�����ٳ�xQ���(8��Sx9���e���֖2�y���g�ԝ�SD�'�SX��j���a,�M��g���$�7m�͗:;��)��p�\��!�,�O�/7H�l�H��!�ʿ�]��ɀ�^-�!�0�_�zn*���~��W].���V�3�TD bFo�׻��E����*��6e&��Y��f+%�����a���%2X�X�1#E9�f۬��Z���v@�.�7_���vn�mk���CqH�Owc<)��|9
�� iD��>\��$���s�4�YQ�k�lF��*G��h�z�q��:Ɗ��HhJi��{���T����nn�h�|��S�=R���W��0@�7���[�G��uT��f.zR�b�T��~���Ӳ�� ��ʵ�`Z�^�֯�>�Gx�䆬~٫8>�\,�2~�R�Yn�:r#�Lt���E�Ɖ��5t_� �v����B�m|f�t�1��Þ 	���^H;�>��ߧ�V���MHVJ�8���ڙZj�4WE�>�R�����`#g��1a��g��>ܱ�4ϝ���l6 Tq��C ��MFl�<���&k�Y�������ܕl����ѣz����Zi�|4�D����FA�);�k���-�CӨ�S�#��ʠ�6Y/����#����$�jif<`����ԴvDq~⽙5Bq�c����h���k4�?��+�jL��D��K���LNn�D��ʫ d`�d���9����ʡ�1����!�g�:��RԔ���?^�}$#�:CC/zB�f>�~$�y#�p���^ԓ^Z����h)#�Ї��JK�Su�~�+��M"�����0����'ټ<�.�χ���>?���J��<�
�
J��	;�`v����N�!��;20Ѽ��F�����,��؀&�UW��\&���|\Y���%ʥ܆��vV���.4Z^+1��k���T;�U�A����8|h����a�:�i<�+�@c�u���d\���k����-�l�ߍL>=pg��{J�5]��H�Q���ѫ�!�e��\GfE��6���+�ۋh�T"�i<$>�d�n.���F�� n�gZJ�k�&�!&��d��4�K�֋^)��W�Ѽ�kؠD�"J�ş�8�g�J��
\�"��DU��(��g��P���"�%��1J`����[k��qs�N^9�jɑ��³B�R�b�}����>��v.[��Q�a�_hX�^pڤ�m^�$�����F�-�+!����w��$͢�V�k����p�L&��N:HL�=�q8��X��28��Y.�)����	N�z�I��+r�ޖ�t�yw^ �r9�q�E�'0ҹ�Su��� �ZC�D�ָp��N�5oQ��G�F��`K �bO�ޣx;�CŽ?��O��q$!$��4���	��,nJr:�Ah0j5���z�{b�r���;�	
�l�<%"+��N|O��EB���� 0��UB�y��i"n��X^�C���̣�b�M֭7/�q��=d�v�$����T�����_��$� ���a�-��Ar
����8�a�Gb���f2 V[?]s�����ݢŋ@�I1C1��3�����r0m۽�.I��BŤ!M�d \U�&�][�L���:�s_/	�=�6Wx�C@vm�����6�*t�5�!�?+|�(�U�w��}�i�_���)�U�p/��*�J���zqHpI�Ҟi������3h7d����N8������@0��+�f�?�![[!���r�J�����Q;�������x�fY��0Ϯ�t�����Q�5���tm�bm0_��c��\��?��jEg�+��Zm	��L���u�I���������V�b��",S:�ch��l�o9����T�\�(�X@g��+���b`*�v�i`�k/����.��D�[�Z����P>��Pgh@r	k��5�[�_������$p���m�*( ڸ-JύCμ�Rp��\�<�SS��ݒ�>���Ec'x�������'��
���4��8���@��ƕmS)�݁�Wx��:.EMИ�ex��\�ڗ��i}��:m�2I��/���7|�R�S�=#�s:i�M���4�媀������m�+c���6�=ռ���W~*)�qH���I�n��a�c���"g��*7�*s۾֫�<%��?�1T��'4���VR�D�F����AU����:t�D�S����e�?�Y��D곚��\�}�oa�G�h�;n�Lj�z��q��݋�FWn�����_��~٤�A�Uם�v��h��L�sx��d�����m��m��vD�ļݭ��UQ�cZTr��U���mO��ӵ�����1 d���ZM�,���~�K�0�����e��g��ST�(Jt#X��'Ke�	d^7�;8^�߿�Ƹ��5�]Ei� �I��fH��u[�{Z�T6|;�g�v�h�m�� �p�P(�-����*'l�c���Ȑ���:_�X�N���	���p�-����8D�V9��kW��	K�Z�7���Ĳ���$�������d��M�M�P�����ۺD���{ǀ��o7�5-w�3�$��"�x�+�ic�$K�rY�r'+��D	u�vD����C�U�a��o�����b�4S�g�Hm0.�[r������R�MB-yǪ��=:��*�x����>h9=X���<�	ĆڣF�������M}��m�I��E"��z�4�w�mL>B P�f	3�+�2:^�� ��x$��q�GT�e��䫇7���I�/I��h����AÄq�mq�SR�&�n���4�-�^V^>v��[/���ʈ��7?�hF�{ݝ��AXlxVHYEB    fa00    15b0xB0#I�4��p!n�~ ����0S����<���"x�O*v��Y�"r�XX-t��ˑ苟a���{6�(�V���ō�|�U���l�
0SW���u2��pyc�� ���%9�[�":3t!��l���{�2&E��5�ҦWmANx<�H}������22�����j�^�������25HS�A9�G����0���X�I: �p �:��\����XV�]�:��9FE�E��,L�T,F� N����T���U5x�����cu*��+�OPw�� Пˉ�-���|��X[B�����=�n3��ѩv��x9be��4L;;�;�Yl7.8���vM=�^Y$蛥'T����B�rM�A��C��+99���eÂ�߸ӗ��+�Do�^J�6L�������7ꅿ����^{`lh��k<lm\���t��2�Z)ҢqE���ϕܬ�r�܋�B�o����7u���������m�:�QM�M�P�1*���$�����_F�l�ۂ��(���b:���� �b���m������gf�en�@A��X��+u7@���T$ ���V��/�g��5�M�����2�q�Fm���;�-�h)�
r��>�T8^��v��rI�}��B-c��x���yU{�tg6��I�ۓx:��ߌu�a��{��8-e��'p)���%r�!C�9Kt��{ ښ��.O�85.�TZLD���/�x8��C��Ǔɛwǋ�rM�Rp�|��s�ol0�L�8�]Rb,4p����z&��Ǳ�RVF|#奩��44[��+4�"5�x���o2N뙑z%� ,H?��CK��%O�YJl��V9��n��g^��V�gW����Xx�UF暁U�h�����ӳ>�˫
=��R\U
��\]�1�#GS�`�"�5��OK�i�ɗ�B��m&��?�>d�~�I��~#�x��a�ل��9ħ��M��^@�'�2Ϡ���R���!����M
M�s�j[�-=�r<��_O�rL7DP��Y1սC<�=K��`���_6_i��_���p2F,��ޟ e��3h�+vc�u�h�יG�-Um�s7o�FL�>0�p�è��2/��A9Y׎�!2�$�˶��A��rQ�>R@FG�=��@�X_�	�/�C���WW:��	4�-+��+C�_}P'��(��kB#��*��������mw*Ly=L�M��r2 ��N��_o18��9'�5�}�,'0�= ��s��2ȼ:�*��6>/i��T;|���^(�03'�)I�o�Jå�1O��Z'�X]�rF�m+�\�<�R=�$5O��0p)���$+��9dos>��y�[<J��1���n��x�/���Dl�	i�0��/یC~����T��������@��aV?�������Bgk G�")�����&�B=�܌c���5�F�����X�ҝ�w�DОԶ�B��j�|ïF͑髾?vx~�owa��NВ� Z�~�gA}@�:$���l��I�g_jղmj�ˍHt���	&�c�a:�HK�o�W\��w��b-},?���������L�����z����P��������۔*#�-�����Z��O��3X���m�`���G�5tx������}�u��1*]�+)[,��1��x?�G�;<�����Y��<vF���,
�ђV�a	r3FZ��|aA]�md'���u�-t,����J��u=킸X�r@_Mg�� ���k-[ �C0���h�%z�@�9L�|����	]/ZW<2�~�1���/Ur���Y!��jE�83z��ݧ8gX	6���qu�N;y>�����J��n�4P�P\]�gM����U��կ�K���Vx�=k�Ȯ �p<���߅��F4���%��z�zq��8iT{d�-���g���Kd9M��E^�8"F��p#4e9�p�ZF��+�S�C�F�ܒz�'�"r�J�X���&��{o䊱j�g�6�����.�h+�u���Ƥ���s>H�������ok�rEh8P�wQ!hk#�F�qU����dt��I���taz���!q�A��Qb��Q�Ĥ��#�鬏����P�S��a�p�L��<>���~s�Cl7����4?gtJ���kY"���Qٹ���09R#�_J��?/�E1�Z�O�A��%$^�p,�������u��Ț�m`�)��  ,���0�^���I�Ö#����.:���ΐ~�r� 7�z�B�t�rF�˴}�L�Kmrd!��D���V�jp��zg����*��$�I^�! ��Sx�B���*n4��\�nM0��Hs���~�k<�5[���˺�3OQ��O�*���~�c���y
��O�~��\��k����`Pfō�� �Se�j�h�����?���pIk�fϛ��\>�<�@�ΦJ�v
j�VN��*B�S�Ϡln�C^fƔA�4���Z����*	�e*9���=g�����q�K�S��J��t�6���G�a��mV7��<�y9B6v�9^�t"��'�/-�q,ֱ�.L��������B��䔵p������W@��	r�w���=:��ui̴R �g?E�K�*�%D��S׼&�9�!K%�:��u����X���S����Kw:�ơ�L��')&$O����aoi�q�M�H?x�B)�Tڛ&U?g���]���M�c������m����X�ī�R��}W�ͩ}x-�r��2�����@-`�ˮ����j 4�p���]vq|��^����O}�O$�<�(Y���mm@�߳~�sc&^����HXˠ�u�R�L �6��儂�:zљ�X�w����v�dH��x��jB)[E��",��	-����7V���sa8^�d�qd�]���7�p��l��(��2��߲l}�7�=[Mmwz[("9��Y�0����}����[�t`�l!Y���#����@�jYC�Ȗ{���'��A�bmt?��K�/x�����W�'*���J�5��Ǽ��ni��g 'g=�Lǲ��L��K������&���S��(^��u���/�!� �r�*g�}�-$.��?O�c�������eJ�(�۬�_���g]ELc�����;�[����g9N�r�ʑ�M�G��g!-����n
$bx���e�l�0V��fT_���D��Xt40�ybX����l��I����7z��߬�N�`���K�{Q����������Yi��	���L����u��[�I��_�J�^o�sGF:YNc��51���a{[9�o5�ݡm&�A�`��h�o��`����5��X����@�ݽ
�0�M>ӛ�
>��+i�}��.����j�&,�\.�Ȼ��!�J�b�Q�T+����@[慥S=yA�JY����r K����_���L��HtfP�Af��a����&ɀ����f�{��Px1���ɗ&��5!1p]bȂ�����Ϫ�㺥!�,[�E�n�2\��5�A�R���b� ��������:k�W����+�G���e�`�H4�$�uװ`����}cT��	c怽a�a~?����S�opw��]�W�x�s��-w{ƅb��������q��y�f>������dc`E����eXZ[`Ę������%MLK+b�p�bZ�6(��!g0~� ��=+��n�l~�Ew,��|,���>*�Hd����}�ća�@�s�Ld&V���'�=��N5��e�[3�@8�⅋[�ն��8_�b��	'F��<m'7Y�۶���O���'��(vH�ȃ������9G���\��Bɐ��Tz����R�x�I�48���U�����C���{�P�J�d�.����������ӝ0�{���������_�	+��J������D�`�@XN���ۛ��Ը�MB,m��\=b`x.���>�����C
^;-�?�	ɕK�c�f[��y��ߣx��s;�!]`���	{�d��R�K<]�8����͊��� �����A���μjsW֥����~f�J�u�����'�G��Μ��>�O4І��4����("ɕ������Ʒ�g���j�!ȟ��j<��?���p���aL
�{:�H�Y'b�3�^�Ѩ���?�$�����[��)�<b��틉Xo=B�X~�i�E�gx_N�~ȍ<�
X��A�2�Ʈ> ����u�,5�v色
�_0ge�"S�V����D��ႋ�{���=[���":����I@�o�i�]�������'ʼ��rvtߘ����s�M�i�W�,�B�-b�pf��n���K5
Mf۔��H��o+L�]��kL ����&��P��y�(����˿�*w�d��)����@���Is�B����.5H�5��s���/�J�Cʣ�E� c�`'�f?�Ǖ���߫ l������ʆ��]���'�0�6����Ό�.�T�p��~{-ޞ��\q�]���5 �vKvru�t\�}�gޱ�.�&�9��#�r��nA}����1܍��@��ӻ�P��r��aLr��OYyj�2
��ŋ͈��ľ�hK~�i�d�b�#2�/7I�r��kfd�K���G���	��%K�@Z�Q����U���Zj��g
��50e���N<�@�I�fl"����_F=�o���"8�ӳ6xd�	|�\[oc�;F �����R���𠂄?CO�A~Yl��1H� ~:I�m/��#5h�K��΋�5�i92%���p��d"��X�?B�9'9�W)�JM�usb������"/�������l�/�qܚ{t��SB?�G���vy��z����gڿ_�pUMv|c���gv?"?���\�r��/���5j���Bp(����3X��{�u�G�aa��cnɉ�;�~�����Gځ=8b<"���lI�_B?��7[󕡼ʊ�²���#���B�.�w���yT�9�������4�ܓ��t�4Y;���ГS�ޚ���wЕ�rSX��?u�KJ!|�v�&��Y#�� ��} :�#��=��H#���M0��͎���W�eB僰�{�WG��p�j��A�huFf���@�@�hi�h���tJ��
*UoVi�ۅ��%p�i{��^|���F*Y��4��t���,v$�x+ӻ'�i!8�$Z.1��ɇ"�>��SS�'kgJ��(��Cu�c�Z���*�e=��"�������hU��$,2r���DPj'�2-:"z�����e����8��_�,������:ʫ��2�(���o�k�Ů�EqV��b�ֳjP��p���}�Hs�
�T�]���xmݚR�n'>�RxȶU�~ח�@z)6��	{RQ`��\aM�t�[b߹�D��jx˸�z׋"�)T��[1nwXg�&R��-�13��@�z�
��Izx�+�љ���ew}TMXlxVHYEB    fa00    1600�1�A�ٌD�x*�����@�A�³+٫Z�Z�$��)-�{S�L�9"!���j��%�����G��PF�u���|B�j	�U>���?�3�F�N�zᶻP�J��fWJ׉���f8~@�(�F�A��({�>�o�H#_�hJ��/Z'�|�cD�r���S�� �Vi�bЎ���~��E�Φ���|HmP8�:�g����r�_�MI�0��Uu٥�E����%B�y���pɤ>�[�别5�ʡa����""��dwT�y'�ygA/uvhAK/�<�0���'m����&,���R��LX���4���؁Q`juX�Di�@̌�CuHX� �O�>����K��ٌg�9o��S���>�E ?���=>̜tk/�4�,v�����m��oK�M��eM���j6eBuC��V�Į�\�q�s�"����>Ë)"�tpÆ*�������$
�=��(��T_m b�"����Һ���~���������N�j䷿',5u�`f�޾���Fu��1�q�O��C��	�2�q��{2�2Me��1�򊆨ϔ�t������lD�c�I�_�{��n~I���"j�n���/�W'n؛�-�,ꛦ�v�2�Q s,}6�R���!d�
$=�� l���K�ã����p�Z��"i�c��F]xؘ�����D~Ю,�����F � )�"�Iߏ,��uF�(ƨ�v��R�K��=�0���z忢X��v�tB�V<U�7>�"�fF�������)���#�t��S���^v�
�Px/��rV.s����P�:�*����58B���c��x�'�`6X6�Z��4{�]��\���c���D[Ƽ�IbJ��;FE^�n�IHaX�0�fg��(�����)�e['�H���g��ăq�I,	���#lI�<H�B~��2�ZL �֋-��[DxNhQ+/��s�Ҍ�m!�)�l,�\�H��!�f4�z$��Y�i�f�:�3����B�A��B��K�U{J:������,��(���A1����a�$r�ؖyGFY3�Q��]K=��J�=��z��/i�i�0�>�V����2�à} �p�����L+�i�?�?��c�/��W��b�Nϲ��d���K��k̩ݐC��bk_n�
z�|Q���lej�3�G�A�V�8E��b��9��:�.=�l� �W�E#�7�r>Z�6�2L�w�B��r��%H��^x�Zcs�-`���4�ʳ�}ɡ�a�tA���{*�֍��CcHׁ^s�n^s���Ά�h䣁K�-���Ee�Yu"lކ��@�	���kP����?��ёo�; ;���m��|�g����Q�V�cߔ�	�S�fO��ZUR��^��ꀡ��DF�)�*�G��3BD[OY�~D*iA�''���`[jB&+j!��l�����Z��1��>������r#�B����P5+z�w�(��I7���|y�9pBp�� f0�Z��]��5���_�b�X�<�0��Ir �Cb��M~���P�d����=��� ��tb��]������P=ɉmII�J=�3��o��H���*��Њ�^�+mųe��^�1�����K��u�B�ɥ�,Y飶�Ahj�@�#</1�a�B�p6@��p852��'A�������Pw�~��>��y�������c_�?	����͉�ѡ��f��{����n����k�ȑ
���	(SG�u:��P(q2�=_�W�Q�[����J�?�w4�a2�]B�)VM;�I�3dǒ�Ŵ�8$�|u��=�Q��o��ioGF�W;�\���v�4/}����-[8p�t_2��nt�;V2�sY!E-�ޕ�X�X�­�sr�<PT"���?�u/����GXk߽�{O�Ȩ'�n�ui� �����%#?� �%�_}�lI��N���ү�������g�h�p+���5��vf1}�>*e�O�=�����Sm�,���aT�xr���`�:Q�(R�,��
s�,Eۖʷ6Xo�>����m=+c8�Fw�H�e�/}׵��a��Ц���yi��[�3�dX�U)��h��O�<�	���]�h���?����Y٥��L�ġB��s�R��ނW��%^��a���CF�~w`5������}�#E�N����.3�X\)b��We[V�+T���7�s[�B/�m^�ӺC�4���=�7�����١��5������XU�<gL
�u�����fV~��]>C�Xc�n܉����gّ�-�;�	� y��4e�{<�kq�D6a�=��o5��2Ν��O5'ô�;p���W2���W��qt����h^��������#�/|�Ls�ǻ��P#��%��ڐ�ģ2��6�y���iQB��|���s#��dlWv��*Q�4�W���wH�Q�֏!���!�3�����R�j`����Q�W�#�"�ͭB��9ә�AYw�Rʲ�X�d��˗Q��a�c�a�Ƴ�>td�Da�3��k�eׅ�y�9��kC	y�6�������˂!�2��!�:�`��^<����c�>nV`������8�# ��U�c�@��������H����A��\�M}�٪eJU}��0�5~��<2��->e����<�,�n8�z��ȶ�=����B�A:�E"d�DT�<=��\&�\'2��"`+��z��5��D}�Pg��+C�x�<n�BI��_)��<;�0�s��3=bM|wU�PWm�jJ]|�Ђ[��0���S�ǁ��F�'�>�N��E��9#(w�]�T����9�NP.�����7�r+qݹ]dMb�ض���>'"y�`Ӏ��Yf6醆�+hU@:m�h���/Q�E�A���iTå�D�A] T��1�澺�3
-�璉���e9r���x�#_Ȧ ������)P�h!=�V���	ý�����8�D�b�
<D�?����@�B���eg2 3/�"/:��#�-I�t��6��h�~~�m�ZM��_5{(�i;�a��[��ȓ�'�I�Oތ�Z��yI���,��^r*���v��Ja��֨h�(P$�<�fGg�wi���^�-���f�͋�t-�M/|,1��Q�z�ߓ��ˎ��$3�N�d�ft��	�;dq)";�o!�^�-�߱FV�4���MbvPP�7���VL��������˜!N�}A�:��=����#D)zH iօ�`UNqd�!d�?��͓�%��cc0��'Z�o|ЫQ��)��m}�7]z[q(�z% y��ǋ%t���w���0AE�9G�����1�}���<D�����0l8"�qYNz�z�e=��n��i����fV�2��Lp).��V�d�I�����J[%Kt9�/��{�Mf�T�EK�?��?3�+	ٙ�	�˧���Ⱦ/������$gG����"��I����6�.�]	KTA6���(7��NmY�G�w�Q��'"Yi`.박��P��͐e� D���p�a��j'ȣa�_�d\q��A�ߚ*�?m*�L\kivo��Y��?��4���AR����lC����l��5ó�or���hDƃ�R܆q�mR���w�R��¹u����k	��4��jT�(��L�U�w�Yh%�e�Zz���, �>�jl d>h�*���]����8��ٶc�� �'BB�-��~�n�Dy��C��S�Zkg��H3��+�u
�����7fA:�_��+(���2��S��F�3��)���b�B풭HD���;�"��:�8L��6ՃL��gF���]��l�Sups�e�b��`��*��ηZ�FgN�N+�������@P�8~�_�U���W,?�w���Hi�rL��D�M�x=>�b�k ?�P�������eA��3v]��8Qp�?��7<�Vړ��ZiY�,�g� F�m��i\Z5S(PS���
D�%#ژ��u���X��8�Ǻܪ����y��~(�5��I����|��tѡ�4�װ�a8r�H��W"n�k�Ὰ��B�c��+�r��[�$Yf��o6�9��1{�K���R���y2�P���6�ᢻ��RC�x64)����A�2�$���컮�z;�ɬ@�1��չs� �Ԩ}""�E�3�W�ln���K�Pԧ)��^�(s�u ~#H�%NϞxc㮛�0rU���I?�M�Nt��-`��~���?�'P.PS2��������{(�0x����3I�B�C���EyY���ebP�U6u��K3XҩSȑ�-Ÿ�*pN�g𐟗)����Ay�JҦ�&2c	߽�0Q�X��[�,Òݻ#ÝU��TՌ���b�;��G��` �)�	-ɚ�s1(�}<���P<�	:ZF�{�S���J��\]iĤ�1��*
�W>��W
#͒�d+�o�_0��8��*�;�B�m�C���-\Q^9�ӈ�J��A�P��I�Yx8��I�E��5���i��ێ�I�\�(�, x��$��l��`>ɁgxGdC�>�aS�Ӿ�C���;�4�<�6���Hb�	��#����G����h�l�aq|��+x��(����c��<_�ig�����/셭@��?^;[Zq HœƳA���=M�Ys�@j�/�{���q
{]�Sꗛ�o`}S�Y�Q	x=����»f�7�2D�=���ܠc�:`����#$d)���(@����a^C�Od�Y�ipb�Y.NNF�+�N��k �<��r���:g��Y>R��»��[������x�ǚu�>���#��X}���0(�d�x����,#|Ohʓ�|(������P��p?�O���O�B���h˪��8ΜO��Z&��ZiQ�~�d��ȗ&5[�`����G"6����o�kD����Ƕ��7���Z��n�2������,�� �2�M�p�]�wkny�.���)�s4d��B7D�/��v��a�=���č��q^����Q6E���]�O?�@Xd;k(@4p���[�j��4Pˍ�Ao{c˚{��-#�Q�^4N�_���T.�hQ�d�84�y<�Gt4ϔ��X@���td��~1b�ϴf<.����[��b?J,Џz˵���Sw؆�����_�N��)8��(9�x�L����|�?4�����#�rH�:r*���ĺ͙Q��0H�b`]}w����Z��C��s%�TP9�����-4C�{jq��'��������<��#J�f�F-v #�X]�+�+�ܭ ��(и�t$r��U\E]'��[��V��UL���-@�˾��J�6��}C-�N�T\��g#v��:՗5�8��k�9���CxC�+�I��m{Х��.g	�����U8C~�@�����BY8�)g�˹=ӈ�-{�]z߭[g��fwՈc_�1�\���=��O/ou�ԧ|�x�?K�șdM;���7�W���?��}��gnUoW-5 �}�cQ!q������;�P0���99sA��H/�3�4!��k�)��op�H݃Orc��B
ͦ}�
%%�	<�)06�(�A������|��3��з��v�Ӥ�<q�A0��XlxVHYEB    fa00    1630�٪@�KlI`�O7�mj,��[,�a�:>D��KK��D��������%�>36b�?X!����M��K;N�Ti��,��s���C����k��Z�A�K�$ǂ��o���$4#�_�b&eU�.F2 o�?V�Ju��e�0�-Ch���(<��i��Ñ���4t���T�4�̈́;G㛽V��X�h�o8�ތ���c#G��[.��R��!l;Ê��G]>U�&��Ŝ�,�����B����8HÃ��FU6Ba NZ"e�4�Ў
��w�� �f�����L�7������`�H1�$܅c�~��Bӝ��
D�y#
�z�!_Ҙ��Q*[�4�rRe���u/\J��%�(
�ź���A�];��P ���X׵�O������
c���o�2��\1F؋�7���X���|/ V#�v�BVe�X�AN��8��<ug4x<S�7�Le�S�O��&��\h(�4���B�a�k3����N}<֬����~>�I��׋�-O�>,˳J%ۣ��G�M=a�����U
�����7ȧz7%�}Ԥ�`����cVV���z�(�����(Q����X��{(��"�x���P~�n%������}�c������]� �ty���Tc�ʋ��/�CQ�)w������5��	�	(�f7Y���BGt���ْR���^���W�^.���Ϛ���Ѻ*��Z��s'��Yx��#��x�8�]��Сkv"|K�L�BѮ��]u{��sP���K1���"����J��1�Mj�K�	�������CC�<{�N�B._e�ߗ��d��ILMO��s��/��{�&�����!Ru�[�O��1����d*R�]#�Y[���3&խ�染5_;9|�3����n�sRЊoo'VН���h���7���Th1q�,kU�T��VB���mu�W�yI=o��H������|�;�r܀�:�b�|�U��v��"��ۢ�5�/1-޾�!·n����!(����N��������ѭ�GЊ^D�I�GJZh�A���`4�l�`ݣ��Y0�N7�풌�D\�t�5J?���0*U�5� ���g
k��L*��S�?�8g���p�l~�B��B�0��������/Ť��&Az��ISک�z���؞>�9T�5��4F�`/D��L��Tr6%�y覩����E��[>;�.�^sz*!��v��k��N��k�SN"^!�?1;Ŀ=%{�������\}$I�X;G~7�Lp8�� �i WƤ���^ ��DҪ,�#��nx ���Xq?�6��$A��W�Z��W�~�m2��l�F�>O��G*�VWՈ�,�̩���+{n� 0k��>Ӱo"������pٯ��z�)<��ط�
�G���i���ؽ�)m�E�r��L�C�i~�I�l�ל��Lz�ʼt��o�ehFI�>���
��I�'� w@�%z�+�#�B�hb��&Sd$N!�у1��9)W��h��a��H���U�!i�)L�x�����s���ڬf�4��JR~IJ���GJ��>Q쩌���"�iI���-O|
�W�_\����ϩ��Z�M���%�[UJ�?P�/*Q�v˲�C�	�^��K_%Yq2胆�\�j�	��B]��r�yn�K�4��/^�ڦ��TVW7��JJ.f,�>�dJZ�x���F�!�^�vE���t:�z%�؄m�W�-��[� �%7}�<��q�XaR������U���1���ɾ��\�9r6�����0�g�o����Ѫ(�ပ;��2��$�F��q[��u4�ra.͆.��'�t\#ꡳ���X�R(�g�#�<V�-w��U��BDms�5Dr��@�.(���[q*y^�`d&���#c��J��r$�ƑT�����N�.e���8�n���>�H�� �؁EO�8R��)�c�\����P�YJ1,t�S�W�, �Q��:�pªi�,7O�]$� }�{�mw
���-��=��є�$�o\:��w�~��0��QigX��7���)�b�: 3����
�����|4-�U�v�E�Ǜ���=G����H y�C� z��O9�壛x٪�G9�o�1���L��*�'�l���UWs�s��Һ`)6"��
3p9��z���"��&9����
�3�4F?ʢ5�5=��?�b���K���$�� ��KE��p]A���p�&3��lJ��٦��q��6� i���V������G�6��S�-w�R��G\Zl�*޾#��3b+T';�����қ���)�7���%aot�D ?q^-~f����%F�Z����|3M���Cb���ѽ�j�"Q��6T%A�~�&��}6�����V�&N���%����hq$���MUO����v�����fE��"Sr�i���?H�C�LAb
آh��4��FW�E�ڷI	Ca�D���OE���\�Xɞ�.�V۴��|�wM�æ���[ ����Vb6v�����X��v�2?aXZ�N�~~�D�Ѣ��q��n��!������e����W��@���fM!�H��� �H@��$��q�̙�] �q�_�s�Δ�E�'�����}��|g�7��\�����Պx���j�k���f'~�YhK�R������ȸD�*�j-I��JS��r��Q]���P&Pӆ���=_r�),eA��;�{��<�� <RҚ�Q%�(8"��7+k;�\��^0\�""�x3���U&MH������bj@;��u�lÞO-"�e����9��C}8��/ɕB�U�Pj�2�J�S"��
I2�]�N���[b��a�}mg���}�Dca�3G��3��ˆ&�'dj�@��h�v�|s��Dް�ww�q�9D4J�㣦a�@�J�9P=#�;K�U;ҷ�b��Wǒw(��D�����k��a��&t��X4����F놪J�t���:@�\r9|!�	m]���j�sZ+�	����u�#K��L�]�כ�/�P29騗��]��UZ$�r�sd}mVA��$��B�{���D��8����!�"�jN�w���zӥM7��ɴt�	�a�ݸP9
�sE>J���*��!���a�L����cR�Q�@s�}t��GȈj'M���ʹͥ��I|��\��_�o��pzB~�̊�7��bZ��|T�m$�L�8=�Ih(̧����1<w�#`�^���Jv�p0V5?�_�f�:�J �Ǜ�F���	\S)�dqw�����m��ߎ@���1�D{���0�W��x��vC�nPp�!��G��Xh(R��_�("F�?'q������/Q�~x**-�r(锾��iDJM~�\����͹\"�� � ���tM��-�֪��Z01I+!c�"L�ueXx���:;v�W�Pk���K��i��	4�}�&�v�?�6����8��n-;��8~$�" �["�8n�<drr�L{�xʔ�R#t���e��xI9)����$�{����Wt��(�.;zlZV�\�e=� ���2�І�ϭwt�q�f�F
�:�œ�^�N���+gq�(:��ro�g'\�:o�3B7-��e����{�	L��l�c��$����e
˚��ە�߮���5�pׂga�(��G?�N	+�-�e��<C�)z Vn�o����G|����3{�3���V�T����Xr���C�g=a��!Z�2�t�_>���Dˣa;d� ���Lg��N���^qQ�S�!2&MH�Y�xy�P�n�GYRu���ؔ#��s2�5�ۜ��\���O�7�YS|�%��*�H������<|�p�C��z���J���T�2[4��ǎT�$|��cXd�V;�-��vߣVk��\�'�VHs��c�����f�r�F���+-�pW�A㩩��	m_��� 0�����!��Nf�Y�$!쌦W��T7�GvF������C��&�|�/�rF�-��r=���Β�)���ʝ��Ò^�݄k�kɡ83u��s/JQ�F-A~��k�c$�^�V'G0�=C�3755|s�2�k�-U���R��A|����h�vOǗٰ��#�O�X<�iI���c�戭���6���7�<�%��*�*��ԟ�����i}e�d2�@���uI>��<>D9�K;�H`���b��¨�0�'���'3I��9YU�?��_��lGG��"�Y���I �.R)���t����_k�6Ƭ8��i]�IK�-����N勊���7�\V�y���}��ל!5�ZY�R��g=٧�r!!������]���F$B������u��OM��@+RޭI��xg�*`F ���w�������QS���t�d�z��ъɡ#���� 3)M1�E��=���1����T��S��Fyb�n���K���-7�T�`��97� �o)�1-�g���չ/1 g���M8�#�#�m�������ӟu�<�HCd�b	��l��O��p 3��UE,{����͋!�/�'���t>9��dKӔ��'�gIT��]��|Un��>�(�\.ZKvZa��<���È6�+Rłf[�j�>�(��
Z�N�܋���!P_yW��a�L�O!��w\�BID�4�)Y(sPc���U��	��~DT� �1��ɀ;�|	($o׿nj
�CFUm�Ikb���|���9�2�>�T��'a�[�a��z�̈3�3"�L-m�0S��Ո�a��
O"\t�re�����NQ�C����[��`�g���츁m@��M}��0����Jc袤�¢B���Ӯ#^��]_��Ɨ����-�-"�K�C@J��	wG��1O�}z����'���u&}Y@�\�IQ���On�ku���_����4g���Or끙.@yo�ħ�.�J�-7���`K6�pÑ�8o�l��f���#�V��}�Nȴ|#����Z<Es�}�[Mv7
Z�Xܖ�����4c_�3�b�z���Y۬��,����KR��}��A���Rl�f�IB��X��V	(TH��n��G̝1t8ǿ�&9G��_J���C���<~ZDJ��d��1Z�n�Gw���Y�ۮ�x`��f����8�'AP���u6���q/�4Ap�$���d�j�t���)y�a�lG��x�v'zETy�/�������b<�[�p���k���-�_ab���܋�>
�*��;ȏӐ�W�|�����d�1e���j��"����wjG&Z�yG؊!�k2�T���i�o���;T���=��s��T�/�a��*&f+��:�~jő���5m묏^GD�=��`v�2�١V ~
�P��o{%����b [e���6�$�+�����)$�u*���{��wd�aӠ#����fi�z[c���A���(�r�	!�I�!�hS���`���g�c$����妹Z��l�,�;�!rJ��̺�l��"�B;`���8��b��gLv1�'ݾIw����k2F��
�����Tj�9h�^�ޜ�<�OT�G��Wi� u�~�Ρa���t.u�rs���o�t���7��𛺺J���5�<�9X�ŌP����LI���MpC����'R�ڳ�ȤF� 9��� ��(	_C4�m�J���D"O�����DCn���#XlxVHYEB    fa00    1620S��6_qh��-$�n� �a�u��t��	��v03��S�Lf�Ӣ@b��M�fsJP��+�s��,o����z�ǒk>����3M.L���"�E���ԋNШ��1���b���_�%�U#�Eq~�ưOpN��cl�������M��c�Rh3ua�{�d�ɡ[�o��}k�S��>-,[&�Q�hn�$;��6r�ۂ`�/��V���`;`jc$�k�h���<�2��!��\0:�NF'����ംT�/�9�?��=�z$x$eA�99d�o5����-�'�����O�[;���^�����E'F�|�6ގ�f!�38�	Oj�x���ީqS�U��'���ґ��{7t�@��2��*U}���Li��GG��M�Ѷ�38!���6�/����b��P6��Km���E,?���8��䯤k�#}��r��9)j�­{�;�I�^bD�������?�b�Cݕ�G7j�k��>~>�<=H���j)c:����R�Ư�\��+�ۧ'�R�~X�ۗ����-{
nt�A��9伻FI�5-�,��=�L�,k|�
���j{��Ub?����$ePdਦ�3��0�}SY<���yE�v`3pXB���.�Ԋ�r,-��
V�f�� %���s��~��th��V��Pݯ� b�\���e��%����M
�r�.�V����}�0�_�$���Xi�b��ZqjQ�Y4�4�)?@k{k�ʱt�f�Y��I8'=��!�Y�L$���+��8���]r?�ZIրuWg���4d���1��A�&�;J�'��\� p�=s�S���7Y!���B[NÜ��_&�^���՜A*�%���t7
�9�uK \�9�JX�'�)�b� ���-�>L�|��2b���Ք�j��g��l�<T���1���w�T�6.~5���r�U�i޳QUD�l��`F���4I�<�+����4����*_:e۶y�PVkǅ�i�c)-\���P$a��
����_s%#&��������7'mOʶ�W��8��'�����Z\i�@���0
�.[-�ž������J`���3�1~�/��E�?�w������3���/4�/�D5c�T�K�2�Jd��wBeӦƲ�NZ0&5�C���E8����b�8��Dh���ƪ��jΕ��|��ٛ	�
i���1T��vp��} ���g�ٷ�9"�yc"�z�5�KN嶑�s�a
�gQ߳\wX��*Caj��{)����zVu>���H<a-�N�CI�������r�@F���ˁV�Z������ S��Nу�kQ�&�޿`q�P�~��`.ޮ9\㵐�{���6VJ��b��v<fT�=���uU�č�h1�}с(/���Т-T�p��!�$�K<ǋ|L|�: #C�ܪȹ�t�Є�AA�����C�{i�Bm��>�nNQp�>`/�ہ:��f?�	��U.k>�StANbtݣ�*`)�Ơ���t� �4��El��$���̣W��@3��h)�J�$<ey���ƕ^>�ʳ�7O-m���3ۡ��ɐU������t��T�Ѩ�tH��$�UuWZn��p�%�m��V!��ԓ#Y_�=��@̰2ge��z�����ZU�t��b����Ϣ���ר�=���*�p�R��SQolZ�*�[���/+�"����ڙ�җI��j��BrG4����_Z�L��F*��A\i?f �^�j�F*�krVO-!��4�Cg'�q���������'X�&�JAߘ}0\�P���=����	�ղ����,$���2�)(<0�-x�~FfiU���&���l����L'�de8��IQ�(�w�H�\7��L���
������b��p���G�;6�Nޞ������V��,0�eƝ���a-� B�m���}����፣@�@w����VՐ������A6���B}����� ���ԧ`��j��vg���T�ߑn�cڑ�����yYE�r;8a�`��3{'� FU��&(S7R#�r��~��~�co��3y���Q,OC�6�Ix�js�%�d>r�"]d�@X6�xR�x�C=;�@�X.s�`�Y�I�����X��H���[,P!=	c��X3�@	�Δ�p)Y5��ov�!�S��㖑.�-c#_��R��k�&�R
�t7���6��,�(;v����A���m�d�nD����v����u0�wv�Ց�E���b���B40��@ǇE%ǟn<�B�����Ü�#��۶nu��ʨ��1W�i=�hxW�z��� ���[zޓ4䤽��fǻ�;��ס�L���@p-�ilU`q��!�n0�AS��OU[i/R���Qd�G��)!l9i�LɊ�
ǩ�1i1�a��4�{*|�b�|�v��<���~�����&I�E���2��W?߁8��뷋x"si_�/-�Q���`1���@%`ő��д^��LcJ��,��&��^w��/�:8���Êʖ���%j�tNӺǴX����ڻe/%XZ�*�?r�Z)���MV�.�)§���F�e�=����iAJ���f��'5=LoD���pj_C��*R��t�`�n�����%i��Y�@��c_�ص�'a% �X��k!F.,7���I56U����9���!��p�\��)��UVB����X������֤��[O��|� �y.���+�s�8QU�Ġt�%б]#�ӷ�Z3����r�
y�LCa��q�ð�s�GHH�BY�x���\�Rt}F+F��w���S����$ gۺ���4��ނwp9ng�>�op�6���9r ��Ѿ ���p!˩��:�n������n�aXC'D�|��!Y�J�?!K ��L�� p��
rڸ"��X�h�O���.y�Y	Y�3��djY��6>Ai���je��TT#��=.�)���U��׿�J��Y;��!)��>�(w8gr-yi��A��v��/���o`~���#�੥ӯ��JI��XL��˖nK�0)��$��aF�)� ���������cUE븝5;9}M�R�����:��Kwv/6'���{"�}+�R?"��X֗���>N�>��3�tF��y���~�@��uDV�j�y*�+���<��݊<���&�� &q`\���a��G���'GRc�~�-�����1sK�#uw8�h�S?�x$����CH���>a�S&<��r�池0i��p��V��[�D���$m�~x\z5(�I���E�U�͙�vR5���?~F�}�nT�Ñ/Q�aV���q�4�(*�H��ۓK�>�E_v�uŉ��έ�ͮ��E�D�ub����-�9U�-�C�+���Y�R�}���~	�[��C�D�&-��_Z�	s4*�nQ�Wt����w���4K@�ȹ��)�<�[�4�,yȣդȟE�n������	w�LIx|D���מ/�в!�
�'���WG��ze������3%� J�$�w�S��I,F3'Q$ ;I�.����_�>�{2�	g���v�����E�E�-n�wԗ>��m�jԭiS��R��S	������`���SQP4E�&�2��`qIr�d����jZ�<�ϧ�^�+��zy��3@�;A�1n��=wY :��M���WV�4���Ǫ/��<~a'�b_W�՟%o����6p�Dw�H�]�Z����3��Sf��g]$j�+�sT��{���:I}��6�H�9��F"u�����>BeF;�ТL�NQU��u�Uj�J!���U0ad}�5��{��~�X�'$��N{jz;z�L��10�U�ۿ8/�o!ƩXҾ��áo�Fd���x��ocj|(ϯ��q����&�{�J��S,�b�5d����u5�����ъ��HE�g�a,����D�]�K��^�
�y��� �q�tU�:=6���t�����߉��$EF�X��c��zj�!�@�@��%-lBi�5w)m&�
���%Xc�K��4�>�Q!S��1)�ڥG�~~g2j�e��v\������<�+����>(v�O,�Z��]m�AU�"����p\�Ҩ�lx���I�W>|�e5X��w�:,���tP=/-V�|�x+�_n\��[�j�ѹ��d
���%ڢ�}d����a�MF��Lh��־2wT����'�5/\��[]�쬀��0}� ~%.ړ�����	g[Ҍ�:c��G�K����h��31ŧ��ы-~�с��0�[�P	`�f'�c��6`��<��� >�%�!p�	>��⹭"��J7���I�<�?^��1S��.vf�aê���8��tj}9��)����Z�7�ha�	Β�7n܆�����u�{���~�2iR���i2e���'1�*#Dj'�����Q����+_'�����B�7�o=�JҌCh���R�z��t�X<�\VU�φ`����E����YTǃ�b�>�2�&i�k9Ijz��,��hW�O��|��k��:H�O���W'���ͳ�n~̈́�S�z�Ng��@�sᲗ�ov��C�;)��XD�E�ʙ���[&��l�	LY*&��q�eR�����|�)�(id����â��o�y���ԃ_`����xZ5;����`^A���G�׭�>GGN��y�a�_^t���P �=Mn�r]n���j�\g�6N��U�I]K%{y'VJ�<�T!�B^�z>a���V�F�:�+^/���=�Y�)��P~/-�M.�!�Fg��rj��}��L5I�O���Q���_	ۄ&>U��=z;�����J:$���$e9ԛt㬕�����y�w�z�g���_������x;A/j"ECY3��t�/��*�P��/�i�i$M�f���!6�b�d�nt2�揰�т����m��<�U�\;��}�w� 1f�A��y��}w�1�!wɯZoX!�� �G�1�wz1^`s�s�eº����hzI;��}`�`e����O6յ�e���O��:��1#�;�$�����q��8w��~(%��gc�y$?��w�^����͍���/K�u��f|OHf<�LQ� �~M���t�͏�5�����q�<����z��e��9�vcei�����[3��_pʏuXm�Z(���r0I�@)�6�Kd���EO����х�*���>l$w���?�E3�� 	a���(ռN��Sd�f�jA�Nh�n�j�N Tq�J�h����g��Keb��"���I<���SH��-�~�w-ʽ\��`j����?`I�Le�t_�崲�����kq?ڿU	�K��'G܈E��9$Oi�B�_3��M>��LЬ&s���L^JԌcLP[P^�~JlJ�ms|υ�tr'|���w���r%�*�7�(��}7����,I�g2e"|�����9i)w!�kڃK�c�3рo�b�b�Ǿ!�F����B���;^�`<%ص�!3��È����[W�PL��d�(�y�m,d=�y��L�᯦�K�5)(��Ru1�<�âd����%�/�5��Ih���G�$�V��(4U�v����լ:8���0]�����@����q��̈́��A��Sb�o�/�%^XlxVHYEB    fa00    1630�lNxj�=�����D�-L`�G���R� � ��>���s �<�5>����~�t��J'��H�	�I]��.�l��T̷z�u�{a,�$9�|��x�L��cx^��kAO/�������Aq�A��J~f��.[�d�tT�w��ͳ��PЉ+�O��U���Z�b;��Ķ��j\r�[~�[�ÛԈ@����T잉(� 
���f]gTD(�م�=�����3~�{�6���1�ĳ�L��?�$�;5?�ۇ�?�	�8ܸG�h�4�B"��.��*qy12tN�q@�j-1�#�V]8�lºF
�E-���ūX��[aM��X�9��5z��GZ2m���)x����{9@�\y�x�|Ԅ���I;��v$F�Y/����J���r����5�υ�<y����;4tbHd�U��eg�����0��ԓ�h�A]a�8�����Q_�t0��Wz�s��q��m�!d8|[]�����;��L��F�vBp�rZq;�?�Y�R�%@��+�R=d�1׿:#��@$�f s��#����1���&(V���V$E�oH�x��I�e��@oI����6�f*(*�	㜳>ʟ9�)˂=��eP�������oM�:.�U,z/wz'�7}-Tr���lC���3��=sK� G�=��'`�x`��� *sg��Yj�%τ5��4�h%:>b��!�	3g\�@d6�x_9��	~A��6�2_�KҸ�e�F3EIP��vTx��=��}��둢�o,���NW
l��`���T0���&D�R��;.��Qwz�J@�'-1u�1��=�$�}�&�#������qS��F��B���0�_؃�,�v�p��!j�N) ��hR��fcnx��cl�)9B'��?��A7	iز��,����><�L=v�Ĩ���R�k��Y,�5�b ܊��ج9ӃZ��S�e:���݈����>���.`�?�~ �|���+��x~^��(:V�G�3��&����2i�\��?�T^E`s[��'�/�a�'`����Uа��u=��-_ہS�VZ���m��d�MK��E�O�6r1i�]��UJNn�'���GZHy�EقآxN�l�Y:�.[{�?8��:I�a
6�҆*�n�� ���>h�V�}��x�m[t۝0ZN-I����J�T�FG?�v�A��"Rych [?��Ag�i�i����Xiy�R��<�ZU1�R�y�2���|�0�:W���Q�z󲂾�KGL�
W�}��1.e��pa�U�8!P%�n�#S��:w`��#�Ļl"�\����o)^tJ�[����E��-iڕ��>k��͓���pbb����>d:O�� jp�[u�d�JY�k���(�;o�� ZU>�Z��t/!(��(x�w�_s%�$A�Q�(��j˴O_hQ]��S��g����em���} "5� �Y��T�T�%��ؔ�(b�kzQYA�	��3�GUj���,���iy��Y�_��4��R�pH�����v�'���u6��9��](�b��!eRE��bs+,�d����k�Gu��_4:�)%��� �1,D9�vB�L�W�0�@~�G����l�r�te�H1ˉ��O=��������i40˧ Pa�j�^M��(V�"y�VUEc�x�g�]�z�&�@:ȵCu�:��&X~� :hkxp�����~���x4{n�ݙ2�1��Q�k{`�/���M\��5|�M�׳]:��8��{�E��wT,C�S��@��Y9�!�{"p-\ة,&"T�=�M[��y5ӏl�I_�,5D8�K�]7��֘��z��)�1�-E�&�����%-
����>5��c�*�ưaI�����{�z��;��B]��hi��������^9�<��������;��w>�F � 3��C��.�Y�� 
lA�7.������ZJ}�d1H�w���Ze?� xωNS�A��<��e���9�^�Ib��Ze�7��� )n�\��0Y!�j;��Fjn0ץ��?�frφ9���
�]w?b���;2*�M�+��SZ"rݺ��td8���õ������Efp��nE�7�ƹϽX�Bh�ZL4w:	bL`��O�ia����H�V���*kyYGcdo��(���� ��)�8ED����B_�K�Tв*��jk�&�Q��n�wUV,��p�Dn�m�ٵ��O���~���ښ|)���G�I?{W�ڴ�\h�����|�X��'���i	�W-���4I�~���������X�޵溺H���Im't�zۻ��+������>� ��`Xdl��Z���I�Jg��YM±���)�i�B�و�yV�uo <1���`�k�O*�g�A�\$>я"h�^}1�i��B7�+?�X�[}h�98}�����\���}��t��a������?}+������dǩ~塀ʔ�Uz�X'�}!�p��5�0��-��q��`��"�4�U���9��`����5z��Y4ea�΢0)օ�� �tUb�vGu"�;����d���R�:���ǧƚ�,�2���D��9ͅ Iv���k�*^r�<�p㙷<�IY�tr �(����*K�x�M�k����S���ǳ9�A�Q�gxx��{�%���W�eA�F ��Ҵ�.��5-ً���Y�i��b/U��潤y��0}9Q��˖-톟�@L"_"t�7̇��ۀG��
c�Ap�F�"m��Z�H�;���~�DSG���	�N̨3r�`����85�d���Tն�p���<2����6�~�;pot�vL�ik�|�?�Dh�Qh�T�9b�r\ޡ6r��n�QH�,|�dt�I�آIi�]��,��̄3�C����)�5c[��~#;N���\?9 �a�d<�����N7k(?��7�c3q@���P������٠շ��W��qC9��~��8�H
�$ ��2i�xv�|����㪹�`_9_U]�^��	����ק��̮(�P@@x���Q�C���XC��?�K%V\	�6�jy����D!�H+�l�`oȒR;e�k��您��̊6��6(�)(�	p�J��&~��\��_0k~c��D�'D;x+h<��}�v��XT�>{��G�Rә$=��!|����C7��YU��F����2��{�� ��C�dP,����D�-X:���:F���"'/  ڰ�yv�WH�.9�����`��W��܂��,��9eF��Ֆ��{�R#�u��?�@z'��aPT���HM��MU.��G�mHL����	��#�A�N3��Xq)-�R琌�s.�g�69��t�Y�� BP���ܯ���nz|��K�x}�I̵��xG9>�ص2o.�8����~�K'y(�ς)+E�V�aGw6���@⟹���1f��әX�:��׿U��}���x�ų苄
� ���U���wΠ�򙕛=�r�(:���#��x��0待�R�0��f�4����%?щ���T����V�5P���yl>�i�)��n�{+A<�b^Y����Hр�ݴ�b�aq��wR�{��(.fpm,s}��d���?����_p��x�>Nx���i� g糠fR�J4%�dA�ك���,�j�(�MQ���*�p9Q�2;*��Z��@�1�gIC,���ⴍ�]���A��e��Gb�;"�����y��ԙ*���p�o��4�9��	�%���G��3@���B�bN�O ��*�ZR�,�n�{���9�B�:Z[�o8��7��l�69f��xQN��ߋG�΂y��a�;�I�m�>Ц��@�4xj��Ij�E���"5��9�-��ݼ=��W�';B�yD|�88���VߟU��U#����t佺�^i�����<�z��+n]r�u��Q�f2�㛋���*>g���9X@;r�������~��c��l�_=t��ۙ���dE򉬥��mǻ'�Cf�=s�Dշ �WAOrJ���Ĭ�Z�f0n�H�G�OU�f~�E�9��v���F��K��W�x��x����:kT���O_L�/#i^Le����';����+_v2��0��-l��
֠�4?�t��Ü�4z"�X����B�`�g�Fǫ$� ֽ
'�C���g���4��NI-�U���%:�.���e�Ȭ����Fy�2��Uד����Q��gx}���dB�-�M�"h��8!���2��TK!�"�<���x�U�qܹ �[+1	�����uTD��o7�C7�dKF7
�n2�9��"�l���ޑ�w�fĘ��#�N��B�VI��x$��83]ז0�>VH`a)@tU�!\F�)�Վ��3̐��}�����J�(MY��8G-S{��-��p��;�$����$U�2�i����6��ڈ�h�K��T(����4��e�x)ݱ:���q��`������+_*�`�U���@�%�'�|�
Wܨb�ɇHĥ��o�=z��4Ǔ^�b^Y���(Ԗ3c�][~��e�L�<�udl�/.��?�t��v�83-(��o,�<ap,�b�@�m��H��J��/Q�
��8�9ȇ�fˌ�8�h�z�$��6%�oZ���g�}�o= ���	�Dc�qY<�6�|c�o9�X�0���o�ܽ���J�Y�c--�Sc�*`��ŋD&�3(��%�Ǥf	�9��^}B�p��b������5�g���ĢҭWs,Y�W�0�ɘ�������~2�O��Gt�X,(M�����X��F����B_�gs��W�SE�[���Z�?��	�	r3��Jႀ��A�9Lx��f��6����,�ƒ(�:�,�+�7�vK<AĴ����@|�)V�7���*Y
R���5� ���l{��p9���!i���f��D�/)\\�w�gw����su
�)e��xNTO��Viזyij���h�l�w�T�X��o1�}zv��J��Lm�WK���V�b�������2��6G��H.��v*��uA�lɆi)�J�A��5��ے!��r�T�,6�iO��m�\��e��kNP�i�Ӿ��w�p��5,�xfJT�`�)7�5��׀�d,����/�����{Ûe�����0JL�  U�r�7�DK\��ڿѨ�xw��<y,!�!:L#Me'_�ͰN5�=�F��V��]y��^����S:8*��^�n��*'�1I���y�S�)�
j񰄘JAwϓ5ME�m����"5n�Z/��O� >`mA�l�!|�&\�d�i/R����.s��}�wq�s�8��6�淵�,H��9�a����7*��:�,o�ېr����9�P�l�t
�TS1H�{��pm����ΡY?���
XKs5m���RWֹ�ڮ�������/(�~��8%9ގ���P�n�
��>H90���l9-��rw-n�=�wd97�Oz�O��ȭ�V��*.2�K�
�@-��YW3���(��>�b�AĊb5�b%�ej���鸳��35s~~�ј�2�}v�"���'���������LM������}���[����#�V��ߧs�!#�u�э�y�w? �-�3�{��XlxVHYEB    5a90     850U��^|�����
�z�`�����X��@G1��(�r�_P��{�5� P=">^�J]������ޤt	��Z;�Sd&n+��f����;>���#���і�(ŷ�Ǐ�T��<�;M;��qa}9�~���B�q��/�^�t��,��o�*���p�!I��J3�2~�զ+��J������V���9��F�W�4g�����&����!4�tZe.Wt��O4ci��M�P��]!�YK~��P�e�U�9���,�����?-�V�m�*˵�Bj�ںR����R��ϓ�ԘW[��o�.���z��ù�R?�s\��,)~,^��]i�ٿK�mNtW��R��SA5�?�Q�WM7�����k�N�{��^u��d��BB�k�&D@����-!W!��i���	of���	͹���"�[ؒ������:�8��WfI�qD�"��C�/%8�r��zÿ���u�T[��[��U�`��F����"q�\W1����l���9��v�j�!xǭ�g3M9\��}����_F�$Xﻪ�lU�ҥ�D+&�D���"W[�V?�A�6tEarBci��A���{r���6H5�,[Y�z-�2���,�db�����)g!���Q~��E��i�X��!���2~Ro]-	K)��@70�<w��bə̿K+�,Sb5鱿Kb$�35ɪ�\�"�n�0S$"���]P̐��(o?@�d��%n�c':�)=�&���h	�.�� �P}"�X�k�lo�XSv�'��0`�}����"$^l�@W���SNbbJ�����uh��`*.}����8B���$��m���?I�&(Q���W���\� �N�؟�]m&���C�>~6�G3�-����MV#�T�
C��V�W��n��D��a�.�����y3H�~jD�H� K��T���c�����[f��$Ux����Զ����EXfOf�U���*��qXL��g0����G �Wq�6<�r�u?y��a���T`�K��ȿ�����?�.��5�$9D@Q�<�O�Y��F��Ƽ4\;q�/����1�.��ែez��M �bӤ.;2O�H�I8��OӀVſ}��ԩR܄d�4���Cq��[���ZU��S貨Iւ�P����?CX"]m���Z%.��5�ey��uMM�<��1�Tp"�{�,��rP+Z�L�`{��@vt�х�,�/�C�Z*�4�L/�Ru��������[��:�f>m�}-*<�F�<��/�t�ʣdę/+����9�pEcu'�K�^�1nI��\l�m�� ��閩2�[��ܒD	�7�*�~��O�x�y�f�i�>%�O[�"�>㛬;Q>�� �~ѰM�\/�U49�B"�Ԛ�
�L{ؾ�B\���������@��Olm��Av�|ͺvYn�܏!��77/
{Vw��䝝���r�e�5�ހ�<Y8H�Y��&4e����uӆ��)�7������C�ds��q0�&����0ܻT��be�+v��9s�<랚F�ΰ!�4y�u�1q���^�v/�8V��:w:FUO0����L�-4��,lL�C��}M-T�AB�� �֣�G��g����x�f}d����#���ei�ҥ �`��Mm9�a#d�����$~7�v�Ȟ�+�C��u�6��� ��<x�C`Ɓ緣���PS�;�m.~m�;Uj��pK�5aP�H�g��xyNM0l��~T�_KWa�)���vM2Y������PƦ��q�k��%�/�����*ͪ	;��g���u8Y�Ԑʿ���^-Z�Wގ�G�v�����uE����_�<����=�����9jÌ�0�TQ'�a��(y wI�q�N?B6�~�6�i?�����$�_��'Uڍ�Ć�'PI�gB�6�� V�a�lQ4�!��>�aֵ�ثnM�!Y9���c �=gPz�^*�M(�-h�s���U�h�L���a�,�T�.m}2�!���@�u3���5�@��L����a��dM�>FU�[���f���y[��	f0�iB�E�]V���#����EZ���o�Fƽ25��)������7?ыO�鵎^@�u�&�iU�+`�i�JS=%%�Zz