XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�Ԭ����gXUr������wY�0�(l7�! c�����p��y*��')��^Q��'P-6e/����p����Ogk���g(��	H�_ĩE���!��.�C��k�_'^oJ�=���Ϳ��]��w�q(N�&xs����[����=��5{@�Y�ɏ�#���<�w�a�d�<�D��M��z�o�"�ޅ�W�~��Sʹ6߾�]�A��Z|���PMI��L����Y�$}
F��}��CZB3V[Eh�AF_(��s	�B�� R�E'�yro���;W�'a�xU �������}1J�RC'���:[e�b�UD��	X]D�D*�}E��1��Bqs��P�����t�?ϣ�+��So?a��e�byԠ^�Vh�JȆ$����Ț.5�T�ؑ��@ڏvE`�?щ�V�~���.Op �}_8T{Gf09(�<���'�+5���l�e�Q�d#l�Zf���9p��W�)��:(N�4mp�>�z��F�x�(D�C�������"+b��K%�ga"�����^�J���o�j��1&�#�6[�ӝɃ$��>6�J�v��!=|��h��E,S�v�繆��JE�X�\+=Ԡ�����U(�dA����@ �S�"�z\�݄�S��6�"�j/7�4؇8��DPnµ]��)�U:�����s�/��V���|^`M��P�·�s��,���Ն��]�wJ�Qª�E8��n�ʃy����0��ZMfMZ�h�R�h�ɾ��s���XlxVHYEB    1ee7     570�=�{I��%��\(��ҍ�{>X-3�)�[���j�O������1a1�օ/�<;�u�f|٬�;���ǵ��s�Rխ��'%Ud�B�p>���mr�[ �Fp�(JA�J���hZ	�U�!��D�L�ũ�Z5���F?�Y�T�>���(��{�p6oYNx	�R��W�IC7��Lb��a�}�tj�P��2M�u\pL�R�#�_�+l��o���|���P�
?��-�!Y��P�]N_�!:ࣰz�5B:'�<��u��Cw�;�9���^� b)&���e��&�������)-��J�>\�����|4��Ǧz��f�4D&��{(��[�S>��K���/��%mU�t�W=�4�Ƿ	���bH��0����@�L�r>�=&'ޓ��R�ݐ�C��*�&55E�o���pA��䙟fvr��4���k�?u#,�]�w����4:��p�AI͝�����k��jبi$Z�g�H�����'����8���1�{?�������4��.���v{M�gnB�$⟳��Ӓ���%��'O��;o�Zg��io�i���~3b�yդV˪�/J7@K��)�̩?ʵ�=+�u��ߗq�%�������p?RA׏�X�J�%��'Dm�}�
�x��8��?]��n|:#�]��?��O�����Hd4�hN��+'��1������4��Zho� {�<	��!)e?4�׺6FjH�0�؇�Ɖ��q.Z��Z��7̀*%�N�h���oi�#G����RI�y��T�@wdeǁԦF'�D�hL�|&�>9=�k��Aih��}��+�-A�8�}����� �.͐yL�8d�O��:����+�0�Ę�n�N�QI�aW��������D��P�Rqb�Ђ  ��&6���`�Ἣ���$���C����<�/|'�4�}Bl1��f�-n�����4'e����p5���iJy;r�MOC����\Js�9�n��4��T�����p�E"!�O}�G�I.�[V�8=��]�������F[��Iö�჉O�j�
#������@�K�#:hE�M@�3:�G
��5�3�YQ�Z����oaUκUk8�]���c�@�2%�Ԧ�+�x�r�O'��[��0<�>�G����̆͵j�H������H��R.�G,$?�� ����=��w��>���-i�r�`��0��L؝�}b�W�W���h�&�5�\'e&������W�9-�"�K�/�1ӎ�������k��JWB��+I�-��w+�T��M4p=_
؍��=Vʼ�-�5Uc���|�gDJ��p*�}��(b�w,��(���y�)�hwc����1���=Yn�d�