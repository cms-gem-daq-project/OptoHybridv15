XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����^a}%e���ㆤ�������m�֘�^*��v:91��S?ӭ���b+�������8=y�	�D��tU���N�9�_�KH�ZS��9QF��(8�9�-���}S�Sv��,^��'tv#�5��3;�h$�
]�%6�����V%�pdyܗ��^+,�f�O�Q�v/!�F-.1V�-Iѹ���!@����� X\?��8~T(���*�G�cܰa��9h�FqrZ�~CǼ��_V	?lyC�"�m|U*�r��l����҈�)|z�6C���h� �><6�����]���1@tJpGv�{u�dS�xu~�+y������C�gx"��ȋ~�u
���+w��Թn�ǧi��U>���K�r��wN���������I�+�^`@��ϘC,/w'5\[�S�Jez �F2s6����\J�]����MȞC��?��(�+&M��%aЭQ�"p�H�g�#5�:�fSn��u���J�cˏ�*�$J���1+��+kJ��%�T(,��4u��Bj%���k_�]|Ŭ� ����l#��I^��URK��.�",��I��cG��&FN����Q�e+V�(�:���24�|1s��WMf����0�wIk��RNT�]��E�����h�d̭#��cf�)g��w(�~ꊏ R�.�X��|S�v�lAG��BRQ�������ņA�c�hm��C�b��@�1B����'
���`/"�m�����?76i����E��.�p�
_�ʀJ/E	15XlxVHYEB     935     3e0�f_w�Y�\y��tj��£G��Oբ�C�AȬV7���1�d�*O�Oе��ܷ���	=�~)��H{����8�!�]c�Z�vAc#�/�3�=��Ã����ط�i��V�g��a��Ƞ�W{�ü�d� \
�N��Z�:}
�<�wO�5��>��z�?7�>`�.i��Y�7�P�Q��߀��}��M�,6U�x2l��0�� �iO�="@?1e�7�鴜% ���i�ǩ���a�t�w��YA��F��*�bn�2�LS/xH9���bNz�_A�"���ri�(�ޘ4I-%W�8�Kw�B�q�Ӝ�F �����M�R p3F�J��*�ڦ��=1�Y��Q���ʚ&p�!�d� ��Њ���ڡ��tCj���+�-Wx�K��U��S��Yzľ",���E0�䧺"fKꊗ��]�_JkƵ�}e���JZ!�Y��[x���v�y4�aΠ�	�s��	�=i�g��0��X�O�㘘est���s�%�,5���Y�@(��O���t7IYu���*��#�'��>0��W�\��ϕ*�f��$���^N�S���\��2ꑥ��ǖs4��D�1�g.12tꉟb'"����<��������$C"�{Ax�Uw�*�a��6`�c���{ǝ�ճ���+�c1�;�"�uW�� !��[UW ���-�[���x7�)	ؓ�`O��e;x���3q��,�dp�l3X 9x�)P�/z�9���?��鏔ї�M��6��bV�<��9}�eG��M��K�AM�}S�7Z$�O���'�n���uJM��'�ܸ ���j�2�i���V"	�W�h���q���y,��Kv7����Oz�\�X�$�$��о�Cu�2r�xi�zHK�gu�kH�"�l��m��{��I��V�|\;�QpHذ©KrR$���rr�˭��ו���B*�+=g�񃊷=�6��G7=��?��b�س���&�