XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:R�7��u�0}3T-|[&�Կ����.5A�gj���cLߠ5'��pVPu7�F18�o��� ��C�p������8Ѧ��p�K�Qw��`l)�������q;�qv��>ܣ���q�>+M�K=}�����)ê+�'�0U�a? ��M�d���Ο:��R�v�0���!�����
�~��㑚F��ADޔ�E}�[���fܘ�	�g�\De=�d��S��P|^���>��L]�W�y#�'"�ƂxgYM
���q���"ŹвD���T��Hx��aq�O!+���j�Tz��¦���Ap��3[3'\0��i�����D9ԣW���Lߟ�/̪V"�l3'�:�7i�m��#�.}�B����@6Q;���jP��g���kG4�9�%�`L��q�
���͞�˔HqXJe�c�qr~TE�v"�Z�&\5������h�D���4j*_�l��ӊ#
Nb��(�>�]
I	��F=u��7
������3�rà�]0�L��00]� F��U"�䣮L�j��ӟ�a ��HgW����࡬g�~��;D�]�Rl�K� 6N���Y�N��T4g\{�=����%��_-���Yy	"�Lg����kj�f�a��sK�Y���p,�����쏈{rn���ꢾ_�G@�:�A:?�H�R��yk�I*���z3��^�ײ}2��n��lVCě��h.L���}O��q�o8w�����ZT��B�A���Z�,�]��eX�w�SuH���XlxVHYEB    3c92     910�p]t��yA�%���0
	-vO�;�W	�V��Xʠ�Y�+ĔR�y�{�$ �Ui�ø��K��w�	g��kϕ�.���Oa�29~�fd�I�����#�㉺�FƗL
?���x�]���C��q%Akq���y`$��o�"��!
��p0�v����I����!�U��^�@�27���������՞B�L!��s��)�,3h�GڞV]vop��0p����6ﯥ���D���f�#�2�J.|��l�1���GW���R�q`y�+C�/G�C��Z��z�x��֑oDx�}�?�~�CH(��4�呂L#���r5�4�̜�ô�A�����nT*�U\~Wƃ���kY�o��'�Y7	��}��4&
�"<0&�K��o��R��8�ɲ(T���
W{�(Xk�w��R��_�% ���Q'd�?�A��+�>�n.�y���M�o�=X3����Zn!�Xw�)��z�O���Ȱ�o�@D���j#g��*�`É����
d&�Tq�����"�*�&irr����l�0t��|�v��5���m1��=��[ģ�
�o�/���������h<i1[�<$uq�����W��.ho�I�x0�d�m�Ú5�	�	�+j{�W�i ����Xf¨	�����y�/J���m���g�q�9�z8��pK�;������k�w�c�+�>�~4��qp-��o-Ժ}�4]����(?�-t��N����YB�_hL�" ٿa%H���e`�7'�{)T�Am��Sh����Uz�c�r�E��E8.px}�R-�Xs�!�w���+�綪^�YI��,��)��|Xgyqa	|քg7�R�L������y��~~���bL��2e�Ͳ����ϑ�	;�^��)Vsץ��m���Q�R�X�r�xC0�������	�B����r�b$qC+,�I������J���Lqw� ��OP!�g�t�w��M^����_�Ė�`�Q��+���#�\Wz|0��@b�M��$�����NH�?J�\��DC�;�ӎ)�>�9Չ��l(HZTA�/v�Jq*o(վ`C�}����R�u�I\�O6�[��<�ꡪU�� �G����Fz�2�[������w�d�l���lt��}k���J����Ňf�v��.�G"�}��˼X��Mm�=*�/�&T*��tJ��3�d.W`��i��]�ԭX�cZ���[콡�y"�b�,@{�FD���d����4�C�$'���z��lc��?)���#}�)�K��v=ߥ10I9x�G�n[@Xz��]phFP>(dK_��|:��h�=B�6���y��),ۈ��܃�
�q���}�9�W��H�m��/%�x��;���A�iK�B���hQ����[��`�-�I��pv'�H��3
�ˀ�,��]*8*Zx�ن�ż��H�C��=�e�zE���yv�&�8�l-s����ŉ��������\�x�5;lLשbx!9���Lw�e8_��3�<�Hʾ/�B3��]#qi�:����	�Mo�)��p�F�|�ޘ]��T*JH��j�I�����R�A<��OFq�R�\�j�+k����"Ʊ��5e�'�x�6�q�gBmj;A��S��c @GG�g&�7��^ ����'*P�rͩ�����~�q��� �7^ѻ~o�H�������ļ)#\tg����^��W�/��H�����.0$l�/E�P��U��	1��yV� �J>))uK��gЇR���`|���M+.����T~?K�s��b��~��� �4�)�̪h�)��sz��!�J�wF6�d��E9n�~)�L� 9Z�̥��:ۉP�F]��v#��S|~�c����-YO㻄��/lݗ]�|&���n�m[��(�$�l=C�P�t��]pN�1�2D|~*H��n��̱1���%��~]��C�ˊ������#��-g����c��G��V����=v���I�o��B�͋>>;݈,��k2�MF[A�(�pp�ȗ�DD�L��$dxޑ]殈�u1�����Ƥ摔��:mO."�G��w`���$�,��̴������J;͙'�0�6�� �n�^����LŰ.�4� �\si��=6j�cJ43���9�bj�{G+��UMm�=��r����;�jղi���ɯ0�.[�a��P��h%_�i~	��ћ��"�ά����:$��V��f��C\h0�N�wf~v�R��W����I�SE���0D�쭐d����\x?͵���e���