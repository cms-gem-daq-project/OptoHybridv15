XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`j�a��l�=Z��aE��7ˇ�t�� z=G�k86�R�KY��QO�A�}� z��)be��o�,�3�2�-g�oC��$�fa�l� 
L��;@tu3�����e@!�#��l ���^�ßӼTc��ߜ�;�37�r߭�֨��%����M�9���]�gs1�>T��m˧?q�l�42E�T1 6��ծm1S�Q��p�Ŀ�5�θ���-Y*~e2k���@�ZCڏ���F�-)�s,�c�t2>�ќ�	���/��J4vv'T/qG�e]���Uw
eV��=:!�?�F�	�>g�FЧa��U���9�٠��c��p�>qX͍��Pfk���߈�!����xʂ�1=g+���!Jנt�r]�w�U�K�U��t�)p�x��0��VuH�C=��r��;��2$�&$�٩&޼�V��L��mtxj#�q�j�5Ry�nH�Zf�6�[�Χ�$�"�YZ5���J�:w ��eJf�q4p�#�!S�e߯���>�j^�!�4"b�}U �����9��UC��Icyt$r�|�L^0�\,���Vx寱f��_-�1��¯BJڃi1DY�t!@0�U�����ҭ(��	�(�|���hQ^��#�?(;�0fI�t��ֻtv�n/0�{vK�ؒ�����p��=
ω*���m;�$�� ԕ.jf���P@3Y"L\m�ۥ^���H���B�����M!ƕs��C�����|���p&w��XlxVHYEB    3e51     a10���{�<A��b�����5�Y3.��yy�\0�/�P��JB��|�)5"�a�gB�2+��Jt��,��FOJJ��?�ހ�8�F�����������<��>Д�4"��K�����Zo�����`4�� ͍����8qB.� �D��6�B��� �d��6T���J@��UAm�ó��1��(_���P�-��� L��C�-�����d��=ݞ����Q��9�k:��_��vR_��5�?��j��`�)+!����k o��[����z)��O�<��c� *oo~ß~�rZ��g}��Ku�~=l���_TA��fFJ�h�4a�,�L����<4]�#X�]����b`�*���#������/�1>I�2+j0z)�9(_�k�94d*���M�/Ξ�7!�����
�C�ƣY�i�%9o��o1�!��T�AB{�������N��'^5)������	��^	+Jgn>J��tW1��o���J	�#��x�z� <�s)"�&8� ���A�Z(STͳ����m׽d�pu�4�mrTّ,hB�F�ێ��<���=�BLC<C�kf#����@�Фʻ�<Ռ|α�_r��E�%��0v��'����~�'�dƒj�����p��q}YC�T� �y��I�iL�L�F�d>Z�Ɠ.ץ�Z��*�KIm���������l��w�)�ZjW�N����/I������T&��?r娮;������^��;��t$�#�c�Z�6��jG�N�+���g��X�R���?��+
Q��S*��5�#>Ȩ��K��"�J��0��Mk&�_u�q˃�j�������b;jg+ș~Ĉ��<�b~�휕�Z�.38��2pB�/�B�|5�׶���)�����Ύ]��lf#��`��^BӇ�M=���hOUp���\�b� �d�"`�-�n�X{��r��9����F�|�o�(���m5�����A-nN��9�,r��e�"F�K�)"��Ň�9�r�u�VI�����m����[��Ӿ��iX|�M�x�$Gv�xl��?�>���=��HȄK�=��ѧڎ {o2�-��q���f�4U�5�|�}E'Cc�][�	DQ$~��x�]��A#���*��ʺg�8`����r��Ǹ�l������6O���W�|� 8�M�ԖJ�?���2�1|�s�M5�+]�����dqG�P������Զ�˒`��n��~b}C��h��0��Y��Mҵ��$]
x��_�>�x>����u�3���{ø��]=,t�!����8���5��5p��h���ʾ�E�e˕qE��[�,�ḃ&���܏ T^��� �La #h��9�b��4k`�=A�ʬP��r��		��1	�2�τ���������CtJ��Y1�8⤳����;_��}�Zt��8����x�.[�3�17��h��ʁq���ژO,��}�S�w��!�;C!��lIP����Ω�����H�O�/� |z�,׻X���H�u7]h�֦t9��_�� i�4Qc�l����V9����OıH;]�����X:k$8��l�t���k�ɻ�ֺ3�Cb5/�
��YbHE\`���:�`~^3%����(_.�RrY&�5)L��x�L^���/Q��ǥ�M�����	��ć?r`@�Wt0���J��i�I���DNb��Ѫ�̓�A�����<��nS�U�!�L�g�(EɥM�^�E�����	a���B!m�O��y��"�R��+�;����@�$�I����7j�{�o�V�O�.%0/�8X�P����l���I^��2|��x��,: ��t?��VZ�x����"d�:��$>�Dʌ���ؚt�PZl����	�N)���dה��Qc5�<�ׂ�>�%��PB����W��N�ـw�2q��f��aѳ��9����l`<��X�s�\��]������ͫ�.�ݵ�҄���P?^��@�In������VG �n֯e��~��w7����䅛&���u���Je������#��S�8�0%�v�0J�����40.$��Q�;�r�� ���hw3��=��� �7o��)׳X,��-��5QW�y$�=��K�rؽs?�Ӟ{26�_�:��Ȧ����[,�I��
#.s���r��3|jp4�ߣ�����~^0y�ཫ�^�-~�G����~�se9��%�Mj'�M�A	��3����h�>"� ��Jt�fF�����K;B��9�c�娯�o(%tb�Ԥ�Fi��sQ��i�Ѣ�]bҤ�Q�`M�?�
`<��pWE����f���
X�����~�&K^��"�_�;�W(�)K{��;Z
��%� �W6�<�B�]x���6�ft�7c���1B&(ju� ��j����Ľ)��(7�S�u�,=����ٵ�}�e��'7o8���6���K��iܙ�s�{\=�`�}%�_C�$W}��ք�%���g�����$��L�%8��9 ZJS�i�a�е ��!�e�p��T%���JF���