XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]z)�C�0=� ��}���m>g�����
�Yv�UFш������[!KC���N���e�-������@O㏱1��S|H�=b:>~����W�+�vP�h=�ZZo	�'�L��gU���1�#=��g�ð��8���� �F�_ä�gg������[ޥ�S�6.�X�ӿǆC8��p����qɵNko��}��(p;t&=j�������ry��[7G����G�k�xp6d�q��w{�#��ɯL��G3�,���n���8�������c��>;oA�+m�D{@����U"f����0)P_rzp��G�Kqr�?��ܹ�1��͵�A<	D������!B/l��O�L��E�����wς�)�~� \,�׏���y--�A����l]'�ǲ����&βL�q��X�=��<+�Aq�G][K�� ^ۂ�P� �	�fj�������|���$��d��X��>�Z��U���6G�����7���+r��$�,J{cye��[?�4.�1��Zp�~��^'��3E_s�D��!�*�R_	Ѩ��|�q��`�gW��UM$�'cU鏛2�Z=�fs�
D�h�"Wḻ
l�P.���ɴ^p7����-zJz
T���V���K�i�NZ�r`�q
K��8���`x$��36�Lx�Vp��I�<	�rƄe�|����)����ͨQ�[S�@��C{�AE����]���]a#c�^�.MJ/oqR��&j�Z��y�����^XlxVHYEB    10b5     410C	���r�w��
�:�9#�S��l��i��a>(7*�͗�u�o�D��d���+����m.�T��� ���a@ɿh�D��C%w�Af�2�� ��C�똜�[C����x6Z}�¼�@�e���m�h�7G���e��ۗ��w[��}�~9�ͳ~�T=S�j��P��w����'��X������V��!��@�+��>�G3ɵ����^XΤ�������POo23=fJ`�8nt�p�&^�X���f~��f�G������Z��(�W��*�9�-��{-
�]#̚s>�����mWY���4�sf",��z����r�A��k)bYw3D�2�NG�	��8@�Eub�2J㶋1ó!�o��i���B������+`M�(RD���^���z$B�_ �5�Fq�dř���5&�r�7o���mw�{4�w�:H�2��� ��LQ��{?�����i�9�R���:��c��JA?b#8�6����a��Q�f�
�Q��N�p�/���}ߣ�!P'~i�w7<���o�+O��拡w�~ٓ\�4�֤^C����h����Ow'37���b8�|�h�2}Pп������W��24�G�ğ2z�4�C��ģ��"���N�N�RvR�?�U4�i$Z�$�XO�_�����hU��: >�`�'J�|���3Z	�#`��|5K�e'����+�,JWf� ���䠔�El����r��[b�6*!ʼ8�W�E"~��R�� _\����D�¡Us�+��e�݄��L3�\��ľ�h�Y�C���3t<��w��4�Ju`/�vR�g����p�=J��Ģ��؆DP�R򼏙aˋS���x�]P`�hCY^^4|2������Ԏ�/�tw<�r�[M9��c=�٠(�X�/��j��Ү],��C�x��W�e��])�$��'��1|;����l3�Y!6�h,qc8����z���vF���Yz�~$F�i�ϊ�"����цP�ơ1����N3秂]ui��