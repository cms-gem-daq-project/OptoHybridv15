XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#���.N�u���.9C��k����|��]`��N��;�/a��AS�F;�M$�' #��h���@Dّi�d�a,��h���h+�%ʛ���BV��a����y��Z�A�%�y ��FN��n��^Z�
�!�h=�$����Z���X���a�ھk%B2l�MV�!D?����Fx��x5��t���R����`�u҅F���r��9�Z���oVJ�:,�ȓ����l�Vh3�d��Zy�Ҋ|�ZS�9�m�#�X+�[m�����)���&"��P^2���'w�5��N3 ��>� �@9�źX*{�k�Nφ�s�裭�t*���`�	�/��R�����S���f�����v#%�Ӣ�Q�� �m<G�Q���z7%���]��
Ey9�^]���Ƿ9��ry���=\j�J�)��su�8��`M;RI�W���FU�fLPqш1��]��PE�u��F�8踖����^u�S�Q�l�V_���b"5����&)�U���g�ڑ����d��΅��h�}F��X�~n!���!����Y�S��I��$�t�O�I�>�SoC4�;]�!ň�q:�n�0oG�u��,�]&l#�V�ab�d���2��C,i�I�\�|5�[��@TRsƣ��d+7\?�].b��[�
�	Lٛ_���"̠��h�� $Ԙ���h8��,F�(\@����qb٣��;@%=@W��s��À?J޹��Xi�&L�wp��g@}@�/w��$�5腜}XlxVHYEB    2b30     a30�:O�Y?���f�3d{�|1(E-�<�pc�ة�-�IE3�X�Ҝ�{lQ*���5�w���������㿡�����(�p?����#�]�FpxI�vj����&\�|ޗ>��	��`�Q�ސߣW;�,�in�
����c����K�rJk���o
��nCeI���oj�I�ڐ]嫐%V
K��JK���ٟ�'�W�Ac�rf���X�D�PW�,���8�L����W����^��[Hs�ѓ �&�����4bE`�o��GNS�%�r��>����hd�[7�Y^��p��P���\�0_H�|7rݩe���p��%��Hy$�pA���Ug�����jQ:�\�±Q�5`s�e�~��?�C�\��~�gD�����=��=e.���$V�zI��kӹ �=�#���{F�C��6H�5�;�c�ץ-��*+L�50j�fʨ�.��g�ڿ��2��)%
�:���T��9oDκ:��ݱ@���l��:	DT����L�,E������Bm���bT�8G����^�����I���/�� ���~��)<4�t�� B��^y�1�)+Z�0(<�s��#�d���v�8:b��XL�j~����aڜ8tx�Lf�t�6�Ξ���!Yz:�&^R>�C��#ǚ9|������/lH�אH���Wv��A$'��|*�,OKz���n���#cX�fu��'���Cǳ�N��|����-��ۿ$VfP�a�֞�-R���y�O��w��C�ŗ���u�ϕc�y��[Bf�xo��/>�*8b� աP��^:����!�� d+S����m�7	�d'�Z6)�]���UK�ҁ{�z�
�p �kb�����3��,MO���~��W`�M�� 0��Z$�/c�R���m�:}F�l��$��M���
0�h�qkv��0
7Lg�����5��
ìL���C�z��o�K,�Y2�mM�ڧ�"��f������Z�&G��Ri<L/��vG��*�?#�
�z�����sy����:s��p�En�\ N�"����t�.w��0�#s�Gg��u���x5��8�Kκ��H��7��`E�U$���َP �P���s�t(e����s�@	ϔ�#5��B�J툏���*i���Mk	t��y]<���.g���S��6�� �	��}6��.A?�S�����@13�G�q7�(J��=�&5�Bwׯ﵈�k3��au���/̲T�CT�E�3��������[�>�~��y��j���1�[��wF&��i�������+�q�u��y��!8�S��ƪ�ri�1����[�;�*i�u��,��̼�ڎp�,��Yڮ2!a��R���Ͼ��4/�A܂����;�t����&��TZ�M�w�<�j��W�dE^��`�����da������ಲ�Z�f7zePώw�����{?<�r��{'�s�W�"����.o�0�ߧv�.�������]�yJ� ��ԛ{�����,�*���Ev\� �Rxd(b�,��IJ]�?� Ҭ��Ǐ =�~@^�	�	�����q'���� ]��DW�y.����R?\b�y�@n{��}0*ާ�y,o�
O����!�/]|�� Q�@ǋ�Ƣ������KZTWO��#
��Hcqmfk�&���v`Na���v���-�X�T�����:�f 7ڭ�B�V��p��	}�5��s�`��.GBQ���%�5|������$���$P�����sA	�������T $��m�$�l��KdL8x���lM�E�D�\%ƧO��ʓTb��+Z=���ܓ[�u��{�G���|��RA���L�_Q����S����E��Ayy�>o�j��HR}��`��t���f@���0�ed��dƩg禇oX8�,�YXm�� k2n�%����u�r\=G��n���l�igͧ�*�>�q�&����F�w9ޭ����Բ"m�JxC��	b]j���J�u�':$���|�]�9�s6�L@��pz��1�Ή7R9K�+gV˜[#��%CZ߮e;�H�|�D���H[h��Ftˆ��&����|��u��P�v�7�xj(�|���I?f�y���K3BEY��K�����އ�(m������C��ïP7�"�C|����R~��ʀǵ��J�gqo;_c0ʳ��t�ˉф���#�%O�/ٚ|��J��V���C��UE�
ODr�~���1��qe2Wk{:�8��'�yϥxs�P?�Ci[���%�]Z<�D�����9X8��3��nLCo�1p8�����W��(�6��S�����`Ϭ�Z+�V~8�|�@v�.�_i��(�`�.�ђ <<� �%n����|���c��3;0�3l̕F�\�򾕺�7���J��}� j�ر?V����:lTx�|���v���*#��bti�n�����@��O�@	y�o�M��L�R\r�h�@px��y����6|�iZ��`�W�<�oP^ģ�q��U�M?S��(I�{|��x�0� �G�/�χ������l�3��Ћ8�U��