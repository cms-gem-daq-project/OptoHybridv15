XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\HbO�ᓠCﾇ@B�g��<b���l=C��n�sF��� ��͇m�O�c�BEm0��9&��W�6�%r�ǧ��u��4�������%���J�9�4�g�)cㅃ%xW�V��m�u7���B��lUڄ�C�{\*c���N�b3`�+q�_=��Y>	M�oX�~�Q<�8��? �B��r)�EVl�M;g^݂�m�b�����֥�
.��y�P�ۅ��
S+�$Бc����&�L_�����ߛzh@�zNQ�>��&�3��{�<>{k㬁�p;4����u?+CߩXV#]��f[���!�LJ&é�p.$q]i-I����%�k�>�A�ے���i);��P�%vEp*g�}V����UH8�Ph�q�����٤.ay}���Y�5?u���W+W"Lu�Y�S��'�|� T�5n�l��<rC�n��Fݨ-�t�+�>\��JӒNY��ZВ��p�'Ej8r�ś�m��WS����40PI\Mq����@��<��+[\I�w����9�-6�JFS�K�U��)o��Ұ鞅�ư,3���
1�_����}P{��e[uzcɃ�����뾬ܰ�Ux��)��6Fթ��Ĵ�V�!���y�Dҳ�?�y�1��jn��bRz7n^��?���J�'��0��}�˟_
J�f���@����W(r���4��i2�k=	Gz��\�>�0��oX�g}Z5�*˰��4t���O�mk,�ܸ�S����XlxVHYEB     a4b     370�����Ok��@�.�L�f6��jW"����,�����U�uu���IE�V�u���
ڥ�ս������x�څ[f3
�=��#���۠��R�\Ү|Ȑ�Q���pWKL�(*��À ����r�Z��^��(^������r�Q������MI�, ��~݄��U˭�	9�-���6�}��� ����� ��1�x����w#\��@6Uآ���Z��-:w�Y�7���%�O�^��^ �p�|a�ٱ�о�n�N�8PsJ�׮� ͤKQ�H��)����61!�U��/���h�f���-$���JN��ҠV#kF�����+$Ag�|>?�A���r�F,����2{�{���7�|#��/fr޸z�Ϣ�_1%�<kN�����000��^�ܮ���ӲO��������(�|��C�pP�����^���{��Z?�e�3^�y*6����x�mO�6rM�yZ@
�����Y�}�c��l(`ؔK��p����"�vK�Q`Jy�g�P��8y��$����O�B��@V6�w����&͟8K1T	�iB<Nh/ ��d��Q���:��([�o��&$��]�Ru1��
ǟQ~*��딧�cς��(z,*t����]Od����y)�i�Z����������z��-p/��ۗ�D?L0����t�
$R/�ЕRɔ^F�S�;�����d����< ��%(z��燅�n c�z Ka41J���_u�I�|}�o���j��ط��<��'�>cֱ<E�H�4��S��KƄ��' �O��,�N[�Y?<HN���O�r�B6��(��P����H�O
�;?���px���Q�O�e����� ���tt���Q�$��vAD��+