XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~Ʒ�Ldj�c��d�:��3�ý�r5>bA�z�,(7��&os��h���' V+�&�*1��1F3|��ͳ
�
ʼY����W��:Y��ޜf����P-�
A,�T����0�":�"�`(U��d�@;?��՜ �h���A�/-a�7K���$�j�nb5�������_~�6}�}��D���Gu�� ��[J�	���y��U����%����/*9V��K؁0Z�KU���p�!��R�%Z��Z)���K��Ru|�j�t�N��?Ӎ�l���:4���U)ǅ	H�z	�'H�E"�M|����	��y�^��\ƒ��	Q�?���\�tX5��j*'kR@j�G��V�2�4"�Oڂ�A�3&���8�0h��R���h�#rf�M�P޹V�=B�l:LQ�&Z�%OJ�Y�pXf�3.�'N}�����RE�M�"-�g�n�s
���b���?�w����(�E�g�����)����!R����h��.�dȜeF6%�����lr(�_���J�(W��������kW�O� ������@�z(($�l��aq!|q�n~�'74q@���Q�9TE��a:ek+Oi�"!��.5�"���Ң�y��KF����j���?�5����U��b$��.�j�?���k�O��}��u"�u��.�m��WT[8�Vhq=�o�S����0�lKo�`<��%��
�+o]���v�G�s����F��b����� P����XlxVHYEB    fa00    1a50\���vox��g����a�Q�7����rWQ����n���<�v����԰�`]�Μ�XH�|D{��B�eK|�A<�^Å��U�BL��wsb�OS�e��'n)�.|��Z�����F�Q��\�S�fi'֪I��]���D ~$x 
N5@�۩%u�G����Z��bNF ��c*�pD������s���U"Ӝ�-w����0��37��)���6��#�²R��lwſ|�.���s��tX����K�ˣ���*b���B>ڒ&��H�?���Jd�k�N�c�|͠B@�,d$�huz���Qn_~�'��};�ּ�E�X)��b�6A+b�*��?�����ۂ�^����4vF �@��ݟ��J�"f�57O���?؀ �3	�6x���]�a!�/�8��̥`�9�{zp��b���%��}�$�3�Z6���
�����,�:K*�B;�<�Os����x��s-=摀���lj�9>��/�7-n��3��CFi(6e4W}��fZj����6��9������	`Q%��[s[��8�C�B��Aȝ[JF�T:�|�5�o�AP���2���a��[iJ�W|�t���|'��7�LJ�S{�}7�h�����4%-�X�KfC�3v�Q�9�+��p}>	�򪪴��ԙ�I������L��n*,�Q��W��Z��C���H�@*�Gɯٰr!�=��l�ڌ��%o�"���|���?��/�r��y�������i�����9!��(�p1�fpU��W*q�1��^��O,X����+����a��B����՞N@T{��uqS6��C�a���"��n!6����^r�Cu�. mR0��"Kwכ�5�$�'�������̽��yPJv�4��W�r��=�P��_\�<�p$�l9�K���V�m٢'*�jZ9�f���&���Oa�<|���V!��3����(�q�+3|π�����U%����Զ��#�"�m��i�<�|`��i��<}C�� ok�i�!_ ����� �c&���8���,��̱�)��tEQ���߲��C$3ҭT��3����	�L��!V
�'[��o5��Sm�B������CB3�ʞx`�so|�V�[���c7ʩu
"�5���������'���i�(�:Y��3�_��N����������ᨀJ>3�C^iq`}l��������?��B@;_h�U~����W���*�3���Ϳ��m��i7ţ٫Ƞ�j���H �D�%\�B]�u2�)半"��-�+s=Q����`
�/��-/���2{�h�[�f&���[4�h��H�v�����fG:��j�(�Fȸ��ZפѦ
��xXM������*F�3�9�n��8XT�U9q)��|�'�W�T��RK����w�Xx:q�&䆺�[��^O��`.�s�6c�:. y,�g�y�o5!%�>�3$ъ�_ ڜ��L9OM�U ��=/>��rA)H^�$�}L����xݏ��#�m�%�@��X	\���	9s�t�k���()9f�P����	2���@k\�%�pJ���h�U{`U� ��l␲@�|;+iM�6 �x����mr<P/{fO��o�	�W�nw�<�n�-4?u�� ����㦨�yI�iJ���5�����@��n|O�ܑ��@�k�<C�kX���^AW=��2g��A'�b�f�.� ��f����Ƶ�k��H��J#ױN�i��*��ґb��qf���nI��W\(a�:Ru�p֛�ڄ���}#H6V�v�P�����m<��d�M��
��g�FK�-U]��Z�NXu
`��5|F���Ie�r�z9Bw��7���z��cH�ݓS�n� �ɢ�!ШG��n�t����em�4J^DYy5��m�L�C]� �g�mt��E�}Hvc�����V��~�������A�6�c����i�,�������У�S:B�L����bK8�,��vj�W��T��g*R{�j��z�?��M������܈g�2��E���t�<�������kGN��	��S�]���uʪ��-~&մ�x1�7&�Tb_&�<;`������?)�5�ޥtm���9Į�{�tN��#�����s\�9���uk���Ne���Q�����֎`]@�El	�9ǧ8vukpb�.WQ�7![�Ї����;Mg5H��MU=�����^�ݴ֛%�f쮁�{�̶��)c���A�f7�u����*��P2I&]C���pm��
Ø�S:�˷�$B'��H_�C�*U���� �pzLUI�ڣ�d���&�pY���~ ��������Y���{�T�":>��چT�(��e�lDZ	d��fG�W%A���O\��ήQ�Rmd.^��E8ԉ�*_[a�k�U��������1p��tV]d�~�)�Ԓ�m���&e�|� ���Cܑ�A�]e����.e�C�N!���5�4j�/t��č�<�����:�����Ų9,S��v�'*�W������)��ĈF;�b3�rHf��ʬ�$�)�_MS`���G��ip����h��t���"��2�1�9=kz��_
v��;�ؙ�o���撯���4g��3^��ѥ��6�Q�H��z|t��F5벀����1���2�����D���b���d�ݝtm$ۢ�:6�RP�5��c�W��\���m����uŔUϺ'9��@����0�:P�I�0\:J��^�K����J��Q���wmc�G�I�Ez7k��a��G�km-G��G��+��pP�}|��޿h�fwf�@B���mQf�^^�r���r|�!���L�g�����zPj����M����p��9B��+F�h����[� �\�01����U嚛��O��7ɼ�1��.�OH�97ۮڕ?_؀��(����?܄SA��;3���~[�4u�L%��ycx�9�/8#��Q������{�|�RD���L[b^�����6�ұ�=�/���`Y�̙>H��{h[e�ca�T@�I�~B���8\��v�/��X��[��e��!'l�sp(�&\E�#U$�·�~	����F����_�@�CT묟p|��%Mes��H��P��~.�W�'�������ש�v��+��S�K�m�:g-���!	2�s�����EŞ�v{*�5���r^�魋�s��}���Ñ;ih��9�YuP�if�?�,Z(�ÞF/��c��1ڝoK�=tgt������V��U#�]���+D�������d�E���*��׻P9B|��b��{u����2r��i��8�Er)��?Q�F���l[�tHP��vlY��-P�UO'bz���Fކ(��V������t�l�˸-d}y`�3�M5؈T	��V�{_7�A��U����3�
��*˛��.���L;ȳo��7�_�����q��1zA�~���\݋�"��f�c���vc��Ql<�;#Th��_6+����,�m�K�,��Oh18g��D�J;����sM�z�1�����:G�Sܟ��1oX[=᧦�D֚�N�;o����Q:q)-�+TS�فȩ"���ȏ��X0i?�\G�,&�]Y����<��B�fe�lv,�F�Q��Jc=�M�􌭯�R��x��r�U�lDĥ��4���J��Tg,��c����ʍz`� ��-�1�������|Tn9�"˜�Vi�\���:ఎ�G�[�ii���%'��0A�[t��Oǋ08�����=���p��Be%>�d�<Gm��'��C�#�{-r_�k(�q�a[�5�mB)����>m�D��l�rjnk��)2����A n�5ښA�a���L�L��q�����Z{�&��'x%9��*��vtw���u����gή(,���I���>!X�$��Y���W�{�R�$��;F{�q�/��̡#��w|jq�������I�c:8.W��ė��F+�����LvZ;(�5S�x��;�X ZOt/����rh��W�L���{�ѺPn���/��g��Q��;Y��U_��Q�l�2�;j�(�U��2��fI3JF��`R�0�%Bg.
���ވ3JbsZX��>�=�����64](��W����Ϙ[����1��#�f�.���O��PX�B5�ѓ�ry�i�I�OS��������N$9�>�?9�V�I*^�-gg�(�e��MM;N	Y(س�u/�~���F�� � ��w	�w�%r^*|��+(1�kZV����=8`���7��� �e�����k)tG�+��cFh��X��_bgy��)�gψ�F5�G��g[7:3��+�6'�n�r����ZL��n����]���0��/Zf����!.�����Lj��#}��ó�%f7j������a��4��V�1dPo����2�����Y�\>}<�?�!\��[D���~�.�����R�D�I�� oi&Ԧ��h[�&��{~�,z��_���LS����a��M̩�uH_1\���.EqQ�D�}X��9{��\��7��	��t�К��
	dMP0�^����Ø�mɟ4�߄@�a^7~�>��n�*$��Lѷ���Ke��L=�M����A5��DB��Sƺ1(��1�a�AM��N�1Y�e� ��IO(c�T��
H�����Če��v(n�bx�q��MW#$�L~�4 �`yr:�ՙs��A�}�S��H�� �5R��x�]�N�_Eh8��;��.	h�KnӞ5��US�%�����w<��P�\����R�@�I�Lj�},��V�@���2���,E��LO�;��.߼MB&y�G���|�Y��W�A̹��e& (W��̸�U��,�۽���%�V<�����ͮ m���b��O���]�`_������I�l�m04�[��y!���V���K�֙4�G)����!%���%�y�\^*�y�`�t�V*0	3^/Tz�~�gm�����~�J����u���~��YQ���>��������ܦ�6E\�[L��M��B!P�Jb�B�ի��PP�x§蒵	�c����@y.��<�?�>�f�����8+߶m--�L�*��Q��c�6U��=��?��a��6z
���$Sա}���mg�KD��(�y�+��`~XH�3
uqIu�Ctje��o�!�ץ�Q��%:#!$�n��g(�Q� �K䉑��a%�=�>�q���/�:$)-� ��u��fU�WJ�s`&��Hl�Q���$_�6�ca����`K���ƣ%'�����o,�$�v��*��@02��*Z��^O�b�-�bɨz���p#W���,����O�}�@�Չ̸�1���u��td�}�~�-P,��,m��oe�s73���w�[f1�Sd�{�v�t)1��3mFb8�S�Z�8��G�N���f�ۆ��Y�ع�/#,�$_`3����SE6U����׵���F��R�j�Q,���ʓr��8
��u옸I|ظr&�_K�A�8�fبBv٦���/���$if6~�;�����aQ�����)6I~�S�}��>B��"枳���{0 ;����V�H�YR]��'�ܮ�($1�oR0����餇�i���25�׎0pօ��iq��h������ ��ʽ�j�4�6V�s;<�y*��mW:�0����M_�5&oq�Ʀ��%����[��� og����}����-�;6=�SY~/iYY����#ݎ���'!��೙Ɲ���7������"�_���S�Y�S99>�"a�:"���39Ӱsowz�z���J"h�h;�fw\��7���Ey��Z@?�/�h�e�HR�!rܧ#����� '+��j�(���m'��8��B�:s�>v2�Z�m�����l;��0����2O�ϣ��>��6�s�SD��ԭ�-���m\�@b-E�o�|�#K�.�%g�2-�'�� �Y��0��G[������Z��6����~��v5&J��*C�5�[�wJ��Z_�.�\��	���i�v�G^���-�k��
xP/�[���'�������h����;��+j�%J�'t�(]�B�n��G�1|�b���
7�_�lk��V��t~D�,���\d�}��W����x�_�?�>rh�R�qL |��T���I�DƜ�;zV��PRE���b\-.�e�G�M���L��r7G�^
z�����³R��=�i�$}��l��=\03��eH��8(�~�����P^�T�;G��v�VC6�ol�a�z	$�e/���?/~z��5*��X
)��o��^���|a�+�U�#f��[��JGL�*�bus��F#�3����nPU*2�A�ģ&\Y.���z5t�Ґ�m�je�2���ډ\颧^��*�(͎�ljv6C�^ߍwd�.�GU�K�3u���[.����3�s}�z�RH��ۍう~����N�}����w0R�t�������˖wW7af��-fJlԱ[^GU�G{+Q0U�^m&4]�C���|����r�w�I��2�+�����\<���8[0�war�B2��Ն�k�fC�@����|�WB"^��{c�ذ�XlxVHYEB    a482     f40"ed�px�oQ�ㅫ��	�����Mx��x�9�3�U@���I�����{-�a�Fd�F ���{5a�/#/��q?�F��?b3������'i���Y���U�n7쎛j4���5�fȇ׵9�ؤ"�J(����˘�S��J6��fk=�a���jEح�8��OM�(� :=K,`*� �����O.#@����x�"�ws�QY�e��2$�0A����ALķ�5���8��T���Fl׿B�b������ FɃ�C0��*�TN�pq�`�4}L�`�^_=%��'o�߽�m!/~݈���)��luO���L�����'�c�!9q$j����u�{��_d氞��S̎αK�:�F�k'��J���!�� ��@>!{aw�*�j�@�y;��
�e��	*՟pn�怰���y�J�kJ=����ё��*}�%�'�o�n�,E5,bpOj�r�6�"1J���3�@"؄?��WһfJ3Վ� ���8�}�<���	���'u���r�D�-��A|�^��t�7��=��t�[q��+���|\j��Q�ߜ3ԑ%��<L��Eg;�;�-�k<h��Re�sZ�0�c��z|O����z�T�W-
���Sa�)O������{ֹ�0��Xv�rkŕzb���c8F��d��T��q��6�b�Ch4���c���lä(MŎ���9��;̾mn�n�ʯDy+tT,�*��'a�Gp�w����i<��>�U߂T%�'ؓ]j�*��T���P������؎�ho��Nb�:�Bҗ�*2�z�9#u/�a<t�]_�e�����q�E\�<!b>��W�\a�	1�j�X�����{�8���"�z�⒈I�מz������7�I���H���hШ�SoTſ���.P��=���*��Ͱ�c�y�l�6N����U��-gq�o�Z��H@ 7�ɞKXa��^�8L�s5�w��@.�6Pn�yw;������>��ͦ�IFn+$> XX����FZ�����*��a˲֎�M�n�x<Yʘ�Lhe~ �U-bt���a����cF�㠼ʯp���~�g�m0�Z�%c���K�&H������`0�������x$������?UW����`�S��;�Zz��-ܹ���]h��rPd՜)n���3��,hfџ$Wa��p�/M�����Q�d]J��
]H��:s�����_��g��4�fd�Qp�|Ý�Dbvm:��q�Z���H%ɬ�ͺO6HS0=�]�MU܎��Vf\P�E����O�9�)��ͼg׏Ml���l�$��Q�\#��C$KY�k�H%���a �?Q�D�87�)�z A-to�� f>By��ٳ:<�s��y�мo����usS���"ܺ4����|;�i�C��iN�y ���˱&����{�߽��+�?9�R�;Ɔ�u�<�c�1r��ט�p�K�4T����ϰ%�]d�FG�d��k`�9�9��j�@�	��zD5sc�޹. B3��"mE��}�=�&����7f�e��rk�&7Ltùr����M�K��[
�l T���Gaj^����&�E
����3�1�
���A�����`��R0&����U�n�XVE\��v���=*���cy�9rb
z$s��O��_���m)$�H������Q|�����׌�ae���r��J�9X]�e�9S��ו�Ό�F":G�~I&^��dN1@�W ������qQ�Ij�L��g��t��M��	�%#Q�� 5��Ęb�~(�-� �}���TW�����M6�Z���t�4]��M�$�jL����C�����.*�n���6��S�u��?��IB�[�"w�����Ϙ�ͤL�rI�S�I���i�x��E���}z(�L���iw�Ϡ��<�pd�h�z3���!ĖP~����zٝg�"d1��7'R�$B�e�v0M���D�u�]e�hU�I�_v6�ԁiQ夌I����5f��<�T�v��[�>�k�GxBԲ�}��h���x�0H7t�n��Z��ܘ�WL���Ӽ��Q�f�{�rz�y�xt���t�F&ö[�v�$P����p�F�T�p��i ,w`M���k*�')D[��ᦧZ��G���Y��_�z2@���9 ��z���Y�d-�����b#�Դ�R�lE;����\Vw�����.�u�j��:��2 �^2�]�����Tϊ���&�I�1�B�o�h��P'P�-���ڴ`����jâS���q֗�\�F�Xg�;��cyo}�0����`�	�҃����+{��f�ܲ�si��^;��]ԁc��+�k��g������O�d�-r)ߒJc5D�(̈́�y�[[��Uv}��<w�k�tv�~��1-���E�y�WO�k�F�?�2�x��j�h�������m[�A��J�q4�z=�����X���X�]�Z�$5̑r���[!"�q:���&<Y�)����)�bŏ�c���B���A�B� U3�H�[f8^�`��a�2�O��b}�懇�+��̬ӻ�G���!}��Ǵ�{a��,���S7a�%cJ)գoD�mu�8�L�'Ά(ש����hY�}��PF�I����N`8�����jx&��W�����bC E'�S;�V���O��t砆��[�Ļ�S�ɂ�҇��4�fč?�	�َ�9�uX���M�ց�]���c�\��9����J���HϱUZ����Iu���&��/��o���=r�3)G%H�>�HB��g���^�D!��୚��ϺAZ����}�5T�p� Ȣ���8`���4�62VL*U��IjZX��G��1� �̙4|鍫��@�9��X��Ua������K6=W��!9�����y���&�V�g<�Cj^ۋȁaK��NV�'��u:T� (4�+�0]�;0�(' 1�K�IFJ�b���ى���N51�9���V���K�n	��/l�E2Z������m=~�37V�q4�^LD�O����w��g��2�41e��a�Yh?M _����9���,��1+L2�C!��fU���R��úѽQ��'�FJ�"D��o17�s��������`vn#~[ը�¿�ǹ���R��=[���/�7U����1~B���hoV+�ؐ��ؖ��8���!<�f�OV�A���9�3�1�1�_�x�i�B�sd�B�g��O##^Vyb�DN��Q��B?l���8Am����j��0��w9��?�<5+�p�E&�R����O�jW~3u	{�ZvH�!�C�&�!�`�hu����?�Y��'.Ni��S�˚#u�h(beA	�(�������u������2F�3M!~L�1��������#��K7�E��eJ�_F)gO�{x��E0�y�7�?�@f&��'*��L3%�Y�g�n��X���_�_������Z7C�C�|�kbW����Iબ�F����ٗ��x��r.Mn#. �N�4�OS�ּT��jMj\��5l7h�J �#*F*Z����y�u����9=�#wWXO�,=#µSH���h^7]�	_��Su�4�ށ��+1i�)�*v6��f�n�S���j1���&�g��;r�;�P.	k��B���-�xaje_��
�K��Dq3�Z>��z4�oGu/ �[,��V��04ī�:Q �~5I*|_�F� ��q4eQ_���L�\����*A_x�R�F |J�N�P�VL�(bw�9r���g��h�beNe�����y[�N5My�O~np�e�(-
����n8�˒)]W�	���+s.�
��k����֌���M�0@��6Y<�g�t*��:�C�w%\! �0��7b�J��G	�wN��a&Ϣ,�G�J