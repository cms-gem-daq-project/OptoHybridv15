XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*l�P��m"Ys�z�n����h1j�LG<��竿�\�)A����5
U�]9��j���D܌l�H�ݪ+ȥ#���M�#���J�s��K��E������36�Nwr�9��K}-H1�L�G��<�R��Q���讛|98_�S��/�Eۀ=��-��쪙s	Ib�u	��e�ORz�o7�(9@�[��o�o<Q4ط9��ה ��@�p���E�˶�����:��δ/��r4���3��W6yފ�4ҧKC�q����oa���>�	
b������b�s�d]r�)!���y�IN�
ͨ��1bi�ĿTsc��l����Y��9��S�P"�uC·��.�V�!�� }�g��a!V��D���}�9�3nV�WP�"�=��1A,
��߃�(����x9,U�|���r��c%�2Y�
��z��sI��!ǪA^� ���|7Apen����	#FD����\�
�C$��]w�Kb�쩨�ׅ�8�W�=ڈ���^L\�!�Vb�{�@�~��fC����USPF�����6OB��r%� �'ER.�s���������$�-���JFGIH�7i~ZM8(]��~��R]���;<,B>�˽=��"A>zW�!N}i���R�b��R���F����_�Y-�	��5kM�ٖ�����?AC1�g��m3�Vv�!&P��
<�-�f%�}�NH��s�ѓ�5z����U05b�]wm��}B)�� ��P�M��V3]��1���e�rXlxVHYEB    1d06     5c0�N=���!:3lR�%�0��t�~G;�vM�Sﴥ"�7�V��8���E�W:�$p/��*��F��7W�����_����"�����.Q��޶��"ٺ���t}8��"��f��@Cj��������X���~{��HM�vJ�-|	�V#��7�Fe�@Aׄ�;�W��w��yĳ>���9���'�V�(�a�r������X�fSK]���v��Z�h���4J��ÖSt|�D����Ncv�!)���P��yx�k����R�g�O[7!��wB��By� �+.Vo����J݂Q;KK�TF��;p��P��P\] \��S��Dߍ^����Z� {��z̢���"v��< �O�g�ri�X���⿼��8<��R�)�mt��9�d��9��a?�EiD������$^K���Y�-���/.�AFWWE&�3�T���hD��w[N�j=u9|�[�����ʨԣ�W��t�q'�0 �2����I��~\T�f)�V�������g�z�*���F��d�"��.�&4��Y1t��{}��n�7*���z+8�v��Z�����m+*vg! d���s"�����Z�Or�T�������y�����:@fi�o�a��)�QJ�;��c��L9��q���-!iT��&�<�_`�ê�Ȉ��B����e՞9Pi(�(�`
jQ����^{�7������]�&A�2
�2�ifw�V'⦂11��q�M^vcf��6�O�J.���b���"���8��f�')E����Fs�6h��. �,_fĘ!/ʧ��nߐ�-�������'ΕLr�/�o��IR6o�D�o�*�dp��!폆��v��a���wwf��S��\�pY��D�����_�aW�gq���ac�����r0z��1��8��c��>��M�<�c{[*tM>֐|F�-�l4�-o��
A�8���&h�f��E�)�ې f��D�>iB�v��nm�1繹l-��Q����y�tz�(1:��V'�RN�E�I�ܨ���pl�;7&� �:���Rf�K�7p[�>��+۱MDx,���9��G-�Ds�n�N�̩�t�v_�U��O>	�3ܪK������/�
aOѮU���[�OGp��-�5V�x�Vq������u�,��? ӟY����+�􁆛΅�&��-�%��ŜC����e��BzZB�8{̏\b�54�jA8�GlI���BԖ�I��&!�"�?ǱrY�kl�K�621zM�x��4���ȟ�x@Tl�j-�u�o���Q�{��|��]���ȁ���Gt�ŉ��K����N��R-�LP��jf�D���2����d��6hV�3�D�f�1,��\�S���B�4�	f�J"�&a���峱ԍ�"����dx�8���=�|Z�nf�
9��֥Q}�M6�Fv�)>�J�