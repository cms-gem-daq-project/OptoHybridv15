XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��޽���@����M����J�L�6�2	��hI�q"�2U����`6��[,-����m�����7ގ(���̰��	��Ƨ���< N�y.1�C�u-<3e�w �9y�����sD���O?}UO*^��u6�\�!���u����C{�Jsc"��q��%m��߬�#���o��D3Ii��n\���`�cD���J	9�Z�):�#�F�U����N��%����R��˩�ګ���e���P�!6'���PM��adnd�����يȯH�Fy�i����u��-wuA����IMR���_�ZV~���k�.R�L:��H��Ⱦ��h%zc�-�����px]x�O_^�@�,����]���2PP,?T�2x���C�w��8�П��N�9� s*������y4��?I@���6�� �b��]���G�>�#ݷ&Vc�J��HMl�3���9�N��c�)1��Đ�Ȓc	�*�/\�4��QgH���U���~F��_�N>�K[i]��I｢��aʕ��$�J���c��.nvO�T�G �	<{!eڸ����MK���ƶg���|Y���K��ǅ�.pw2z_�(��Թś�Ņ��_ׂ@�e
���X��=�^]�5���V� �EB�ƈ���W]'��l0?Z���_��k�hI��!�g���U�ᐬ��`
$w������)��O$X��,�TF�}�p�_\���&��Em$,6���P�C�C��5D���uy�q:@��XlxVHYEB    7a0a     c10�/Cl���]��UyZ���q�u��m�6]B���zv��N��&Hҿ�X�Rܵ�� �]m���b������xaQ�������:��s�d�Ie�4�ƚ��P���)SM�qf(�ٹ���
�Vt%}h��(A��/�h �9�/ؗ�r�cT��K����_�����m�������(K���5�Wo>me�]���+*氦8d!LMr�$ڤ9�&\w3u��n��ɈA�t�l;���Ճҥ`A~���fޙ:`����1a�j⳧3_�9;6���x�+5��y���O���s�I?�и?[�IV��d�����I�]0���������IԦ}��B�O{�j��Y�~UU=���4z<��'8T	�����؟M[F�-����E)/�i=�����[0�]��X�Nuk��(r۟�D��(bps�.f��k�g�:�s6>��m% ��Lyqp��z�l[B��f���Q=q��/�F�Mk`�Mփ��aH %�)�Qf��lC��I����c��S�4��I9:�:z);��y�K��I���N��yx[������ǟ��tF��C�ω�h�Wr-�=���6��B���C־A�^C���jz�/�|�ՊF�p7`���Nڕ��
񍬘�<�$�%f�TaŜx��l�}���k��~���LS�J!����2�G�Λ�F������_~T�I@
�g;�s�JdŶ-� �Ɍ3�|�	C��/�c�H˜^T������P���,"`m��[Ө����q�b���S|���ͧ��{��[4K(P˞��T��͢�_(f*��9��"s5C���%�,��^������.=9���ߴݘ[\����Q��]�j�Q=��n"��x�R߭/!�(
��l��YZ��U����&^}1�%���&<5~�,F 1�&�x\R����t)4OX'%��H����<#�7������;�F��`j���*��ɣEv����ipbi_�%�C(��q0���/��}S���iU�1zV���)��}��ؤ�r_X�'�H�M�*�c��x�e!������B�}��\��e�hʈ���c��G���Q�{��2h����V�߄J�g�.�3�4Iq�Zjk�`00u���@(Z�#�vt����M�G���E�����r?�F�OM9հ�.{����M��i��6�T�Jׄޥ�_�D��;���^��߅��r�ȹ������!�#���3 $����z��p��W敢���ɫ.�
jiZ��2�s�)D�."��q�9p�w�b���V�b�?Ŀe��� �1|	"�U�!zÒ"�9R��D��5B}��1qX�1�Y�	%B����&)!��Di}*���	Л57qDA^����V���Z�!s�K_��,Je'���av}�f��.�� ;r�5�p\�E����O���8t���]*�B�uJ�8�W恰L$x�;p���_�e���ey�1� �I��+��Zh��6'�� �Kw~�)�tͫ�)�bVC ~}�Ȥ���C�t�v�[�U���/J�F.��V;�ǚ���N)�6�'��^�C���	��e�YqpCZ�+1t�Rz�{��5{TЧ"���`��f�x�ͩd�q��A��"9XG����5%gv?��5�K�~�Y����^��� ���-�/�!��k��{�R1~����u�\Ȩ='1豙� �rR��nuX
�^�����,�NRa� AW��4�ӽ���z����e^�t�[�������Ȉ��:��6v�c;a1Gc�G٠M�r'�n\�X�H����{�V����U�bhf6��e_u�q{� ���1���5"^%Y!w��;!F��)*c�#����:cd�k�Ҷ��r%��4�2�<d��N�Z��8��>{[��G�^/E=�==����G�hg�{8V� ��i\h�-[�o�JΩ��U�ƕ��h��b,�n��`q���-����>�%�L�����qI�҆t��Zڨ��VZtM�W)]xJ�[�`�b�>���t�Ee��_B��I&�v��J�:�M�yl�Ջ]�n�);�3v0vM��$ڮT��?�s$a�S�a$"���u�����h�5��4*��.��퍂�>�0�3��B�W��(�on�:*N�S%����٥���3I��~����P3#é�ֹu�C �F=TH�Q��}t`<ȃ�s;)�0�(E*�x��H%�J�����080��ꌼ�O��aW��.�ح�B��ȁ�~#L���	�8j@U����`fa���Q��"���Hă8K�\\��u�CB+��7T��_��.���o��/�0���Gyfv3�p�+�6�Q��v+�8j8�h� �C��h����!��{,%i;�E�Z/��ث,+1�w��� ���V�l�]y���E�X�������?A�.J�^�C�-P���U_��㫽i�2���"G$H�ɷ	�oʍ����p���,��nJS�����p�pU�ko]�=xj���4U=��ݮ:te�*��sM����Z;��n-��8��bB>聾\�P�~���Ӡ�_�}MZ�=�J�	4s�I��1��J�d�2���n��M]�J��m��I�D5[M� &��ܼr˕gt�ڿ���QBk�Q`G�«��$[����R��)��%=|ۢ�J�bcG�����gjULZ%���oB���_���f�"��L�BMe����;J�F,=��8�+������֬tM�O8�n7"������Lڒa��v��+�m�:�|��UI��q�!�Y��
)Z��l�>X͉S��*�\�U��E�[�o��d��p�͛����B�
AZ\:�-����c���9ɝ��ʮ�/f��vP���̾ms2A��h�,6ti/�^u��������eu6��@j��a�#Ω ��O�ҧC�{wX�p��5��]W��Pg0g�ŉ|&B��E�B�9]`Ay��{���f��.6�gI�5�^v�[�n
���z@�.k�o^�c��`\E��d��CY�W8X�