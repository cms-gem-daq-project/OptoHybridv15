XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6Kr�A8� �8}���T��Bw��_�PYi'�KA�p��!굹Ù;�����(%N��:g�PM��O� ��~q�h>����4��ҕo�Z&����I;���'G.�سqO�ϯ�HT�C��ʖ�q/0�̹�x(��kD��{\jM���-7+�R�)o+x��F������a���2�r����*�B�����J����Q��	���nǮP6(��I�I
��ٛ�v��4�a5ר�G�����>ze�Zc����?��q��_��h��t��v&<v��{�(�5��p�%�m�Am$�.���d��)�Q��c�#��[!ւ��?�/a������
^� �9�b�G;\�he������g�Gsa�.�:hd��%m�뉕p�� ����|���k
[�݁E��?�:V*���m!��v��
�ĺWs��� _�g:Y�Ή�F�ᤔ�bkp�WdSs�����È�^(��Y�t$-���m��ٹ31�\	�3����-��@��$�������S�nmr��㊃�PʛM/�+7�0���>�x��G�˙��S���<�����g&�a:a7i�|Dj3����1V��uvm�n��!��/���s0���1��֯��0�PfQ�[ ��'�����L2��O��$IkD�s�|��܀$�^4)���n��d�Ē��j:w�KVOv^U^s�zk<�r %|�vzh�k�d�|E�"ޡZ@�vi�;"|т��}p��z�'��1?���Q5�N�	�}%qV�!�ꑡvkC��XlxVHYEB    2fb6     6903��S�DM��1�׸w;=�yD)����_�3JO�,^cm�.�?X�]�E�m
(� ��y��U�
�}��W6������?����#;[����)�.�C�b�h��Vcvs�<F���z�`0x����Vԯ�5�sx��!nd�{��������rF�V���j��k�q�5�@�)J-Jq�kE�-#���P����LVǅ9��2��K�d-�"��롛&F���$^?�D,����� ��s峲0)o>�5��b���`6H�CP�Ae`o8�_��紣;`���2<�}�y%�������k����rt�;ʫKϨI���4H�GRr@�z�t|�z�-��%OsO��T��'*�0��<�qzJ���O��E���1[U��M���jWGP�q��y��6��h����z����v�l�B5&O�����I�y���m�w�2\��
\�jjΙrhR*O��m�@TN��[]��+�[�T�����]`�?�,�����0Sz�[:�uP(:\Q쐾H�>��^Z.�2��f��$��+W9��~�2�iAp�/��?����[���Wi׋��'�ص�p����Gc	L�|��aV���D���?Y�=ZH��"f���R8�[r�\�\���=�;���5�k�Þ���c�;�K�R��̰XV�w�q�y�sy�z� ��Q�w�|�~B}ϕcKj<.WS��[s�gq
]���LD+���8�D�"V���Zk�`����N�]�!���T�C�{@d��-�+[0��avx�������G�,�^�òc=;��ﳪ��!<\svT$թ.�_f������u�rY���	�sФ��\������U����
`%��4d�o�v�a 13i���h,V�;����܂��32L٬�[��Gp;��� ����~�  ~p���E<ԁy.�J�)PQ�6����q�95I:.���X�{���
7�&��՟�AH'�izy(~@Z�q�����a}�Hs�k�Bn@�Ծ�`+>_|������_��#���DU���P�Z.�W�j�� m� p�á�撦���R��W>\v�!BS��������a���z-��r�WGG�벨���yU:�,6	/+w��9	����Զ��� �P�$j��ض~�F��5��9�~EC�-��V@�+hQ�zO�vBн�q�	�d_����e*B\��Hj��߲��vJ��3��)U!��m�����X�r7�C�˔LԺ�}�N�|�����{�;�%�(�P!��%���qA���㹱Y) <M��nH����/tw#��D�.4K�JbΜ%��ü'��c�󰴰�� 	��,Js�ST2������ ��Gj�1��*��uJ�i��h1aا�&QҺ/�>���VBP��̏<���
@����#���@�U �i�e���oq������9���kb��a�hWp��59G�pT�_/�,�-�}���&z
[�=�j@۪��F"�ټgF$�/FPϟ��!��FT�o��5u�������wR5S ���Э���Q����/�����c�����R��`�����ق��w�� ��N�i�4�y�<�%�Mf1�Йڧ	R���M^M�
Y ���:9���4�����S5so�f�