XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����W�[��N��	R�}^��j����SOWM5O���)ܕ$OP���O�N���TR�
�(�}l 9��DVC�9ƛ�o�+��s�17Y���o�����tt�a�m��S�����d
:��(�=v�6��|����ei4�1���CO���G0��p���![`,o�]��4�%�qH��fQx�D{Kǰ�Z�5��g�E�n�y ���L̂-ݦ<*��W�̺��V~������x��Å�R�汛���]l�ʿk�X�X� NόS�/��ƴ����to��v��$���niG��,?Tv���+��<yh��Й��EM�8qo6�����?%I����1=�������h�S��Nv֩Ԭ �)��� �LQ��'o�G���l����%�|*7�K	�s��G���$��`Q��q_�u�qOp��>
�T��.$Bε9>�w,�.���\�h�������z����J��8�&�>iJ���=ȅ���y�̥¼Tvf�)�
Xfԩ�
��-����B��%Yn�6�1�0���F���A����co1����<-��6c�5f���Q����=l�Y��ړ�2䰸����sd�yb��r���r�jjvJz��X�F�!.���"��S������%�r�%g��<���;����Z�)6�����)�3��ǻ60;<�x����[�I �S,I��s����X���lM#��Q0^��?�Ok�ĥR9s�c��HO8n�N~�@S(��4+�څm����94gXlxVHYEB     686     2f0��{�9]+�(�#Oq�Y�yΗm�K�P��2��T�Z D씨����Ȣ��)@��}8ͪ��)�U94úd�܆����^Vʢ�ˢ4�	>��]��%�215����o-�N�����K�˅P��r��t<^D�6�F>��+�����=��L/�ư`�1|1�!�p�^�30�l�ex��Th��KzY̔���Ӏ[�'�4�&���?a7�D����qoVJ�����"A~�$$*X ��v�v��˫�y{$�Z�y{@��I=q��� 佯�;�Qt;��`�Cj>��Oִ��KLc��㩠����k5��o��P����i)��c塷燪�?���e�
�]��b*��t�����/��S�f�TTZ�b
�� *���|���?ptk]z�����w����s+;��լ�MY����#��Ms��>��7���n�ٜ�=�z�����nI�S3g=������R$�/�3���
���6�	D�����]�ia~B)k-�B$�a��E)p������V�'}��L��֭&��> ���X�҃-���P�������ޖx�B��R��}U�O#�oi(M���i����^��qO(��`
�3���J�Nnu��� \�pV�����EM�-[_κsh�`~��vr��
�;ڙ�c\'�����惯���0���LJC���	#8�����%�[�#���J��j�Z�(M�ũ4�jB�9�=���\�iU-����
���D�?�