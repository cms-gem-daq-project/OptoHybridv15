XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�&�/�4�L�cE(�dCqBtz��ɽhE��x<L˸����}�[,r������`�&DoQ��0�wC�#T+ѱ1�x��[)GdN���2�[$�b��N�)�3[ZQs�X���� Y����3��T�|~��M��a���%͌,�]��KΓ; 8@�O#A��&��Ģ��$(���w���ǅ!ԋ&���eS��B�W���,z¸��\�=�:��RuK�l��HVI�:�P��c�����2PP�n��|�o*�:f�9�>�)�#1H�b�-��H��������.���|��7�a�������Y�)���ɹUƞs��r��X7��0\ѤX]wq���T-��:"��`�E՟_1US(ey�IFDP|�1�����B>�
��L��U�ʊg�r��s�����4���VW�,U�Y6����)Ùs�gsWb'aOn�=0�Gj�"hz�U�[���	B`�ڧ'Ԙ�q�x{X ����Z�ͥr�"�ϓdX�����ЩVYr^���5z~>�+�	�8���*H�M��釄�����#mª��B����Bb�LW��G���o��"�T'�,�s�~Ú�h�T����6sXԁpL�Z
~h������;ُ���k+��kDg�����$q�}t�ت��\��6 ;w�����_�.c򢯰U�A��w��D}�F����5���Ή��U�$U ��j9��ۂ^ϊ[Vk�Yg9�X��v-�,�ڑE�#d!�7�zc>�~8�#�Z��FXlxVHYEB    2861     8d0��JX�N]�+��%ek㹬-�W ;넭��L���2�Σ�d���]���WY��:�e%�`��;����Xj\l���grkTm�|�F"2l[�W����W=�@�*�%��-��s���I��`���v��FoF��f��53�-eʉ��<�Qh����f��l$�' ��p�PC�"��-�P-��H��'��a�bKah��:���h�̃Х�a"{��R<W��E����jI�����M�fK��9zu����6��+��T8$�-��bI�Y8�֟YS�GF]r��խ�l���� ��҅����R �:�?�H4�����9�m���7 po���H4�܈�u_�p���+����P��/��xb{�����O���� �Si gϝ
BN?O�;�%^IQ1�I�?)�Vqn�ʝ\`S�eyà09H~��^;)o��3Wx~4�aƞ?�0:	����i%�v$�������#S��Kʖm�����^�}*З�8e�N�^�3��iq�}J-���~*u
�E|�Q��A��z=�5�Ϯh6��w���l@��s��&�[>����>���o����	�h���o��kW�Xu��%��'�E�wPz�%�*Жބk�_ L�5�T�1��9��ؓ��&ѣ&��:q��Z�yhԦ�&��u���~f�ꓣ_�J^�cK*�r=NȖ�}-�SB'�Dy`�~(���7�z�����D�-�z�Ə��:^V��Dx�U��?M�	�^P���~�*<� ���h�W�Lq�)s8�k<�:x�8f�J>��E*��-�dr���I|#1��vMwD^����K����_4�]-	� ��+Ng�;τpj	�u�}��޼�3�'�+��������� ���!�9�pq�b���� dlx~�	YV��z4���^�P���2�琒�:��<ъ*Y͓lO+x�]�'�1���سz�0zn�j�|@r��L�XFIMH0��c��� bD?�wa��fk��/QT�%s߬g�!�q��Y���Ŗ����?R)`*��<�\m�Γ���
|�b;s���$a�ҰFOŇdc�l�-5�E����+�`���зɒrj3.�����Ê7ztug�d�����2�a`�%Ə��Y�S������{��6����Pk�1���	M�+Sݑ*D�fU��t��K-��H*�a�x�l�Vo��O�5�!7�BΗ��/[3C9v�|�A/��d���CJ�5��Vo�<�`+�ޫ�Ճn����Y{V��Z�m��(BD���A��Oow�/����u��u����ң������~-��LgyVbJ4����7�N��ó3��*�wQeJk��o /I\���� 	��{i�N\�H�-]=p�r�(M�T{M��HR����dDP(�h��]f\Q����@���>r�L���I&���b����)��� �4D;����K���[���=Z��C�i+]w�<����h>?"����h�I��VZ����|��~,�;o�q�����jb=�U��}�T�9��)�H�V��D!���<6�8�c�p���~M	#��>����R�PYk�A�uG�/�ı����Y�_����tl�"����f��X�&�?�b�p_F��ŜdD�����NcL1~i��f�k�Kt~�TW��ݫ���Ծ)�E
�~��'u;f�v���ʱ*C\m6��/b��Ei�u�\��8§��l���"bt��\1�?�% 0�f`C��6���;1gN%<c��N�%�2�7s��{z����fu	��v�-�5��hc�s{9�Ǣ[��P"�m��}%k���3b$��7�&L�8�q�y�z-��b�c�F� �w�/q<t�[:)�p]�h����TjX�٘��w��ǻp��/��Y:i��Ćk�ٟ�����W��3������&�'����}�F�jX7�[W�-!E��]�e�K�5��';��/��	
�_`�I8UY�6���)kaEi�L�@������D��װ��M�̿�5��m��Z�s�h���K�@�������-�����_�<�>����A�D���ǰV��W�J]!��@<�l�Gؐb�h-�-g[��zNOӑ��}C���qZ�s�4�xT�M�ـp*r*���ɒ�PI^.%C{�
h������,�nN/*��{�;kU!���z���s�����|���k�k�+�kÞw|�7��s��;�c�S�7�