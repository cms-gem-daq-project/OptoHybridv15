XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e��} ��Δ���J�<yXݾ�(�����"���O4*�X�1R_k��4����S]��V�6��|@Ynbjx��P�{Qꖱ�M�π2�j���@BϿ�Á����xaűh0s1OM�jՠPH�9P,�̸qqz�X��,m"#ɜ7��@�co8�t'w� "�_�8�6�7K�%\qW����^6$���&[�ʝ��Y�Nu�q������W]��x�Yo��=��xSY����m��$��!��m�C��-J6T�N1�}&�ERۻv9�<N�r�y�6�a����R8�H��"RȬ/b���l"P��>=V��]�H�~\"�H>���[ȟ���yuȲ�����;6����U<��5%�G\_P�����IV�ʀ�.�HŽ�t헺j�c�&�!f]le����YU�U<j�3����*Ίت�,&�����M����0�+��ȿ ��n��%�[����޳L��Y��ID��VN3�y�"��k5]n`����{Z�\,�|�(kC�4���N?S����$�	���;�:h'a�Y1��g%[	�M��X���c���u�)����K���ҁ�/P�ۀ�<����Z�\2+�x��@�q�^xO~~Y��r���3�$��hPPh9�H�-����gmI� �Peob&�Y�:���8��"e����a4�bF�h��J����F�.6�Gz.�؞�"?�2@;>�LQ�'F.1��C�hfY��@�۽�����cu�쌊�+�.H2�aT@�:�XlxVHYEB    6faf     c30fM:�`��;���1���������N���<�a��[2��S����ε�ߝi�-���T�d�k�g�%pc!X����L����&�u��� J���>�"d����Z<�}�4e�0:B-�K���R�_�/æ��U���d�"C��H��i̀�����H��%Ip˃9o%'Gm�P-��?h��|l��-5��A���_u_z��;��0���<�e4�A�)`p_4W� ���1���*��Wm�~���2XE S��ᣒ9�	ThtE���\�
ˡ�đ�Q���P�2�����x?,늤gL&�F�E�*�JmL��%�zp8���?Z�#��M�P·@,��qL��+����sb�ӥ׋l����4�ڮ ��ZG��	۱fKx��VS�vQ��L+��1�O��;���J
���d���B��w��~Rts�*(u^��Aم6��6=˷�I4�����7K5r<����K�q�+/ͪ��?[��\n��\�/3�Ou��D����Ë���Y�ĸ���ͨ�A	�ÿ�*зښ������fT"�M���2��qi��>��O�_�v���}��|��56�kA���h�?���+*}i����{����g"P�A*9;�a=�5��F}��Q��|,��9��E����"�� ��b-5���:fw�6V�O�}�)tX�)�Z�(�����u��F	{���ܪS�]��dT�z���)�A�9FòفzyQ㘱+b�+Q4�G��g޴�c~F'o�&���
��ӝ���4?D�+�lH- "ݥY,�M��D���s�nF��+�+s�;�l~Y��V|pY:��3O+���Ak
�n@�ߠ V	���x����M��4�;���Бl?����f/]�4s��m� �*��	�m�@iA��NZ��0%8f9�F�Pyq�?���r���)?"R�G+�}R����ih�e�D�!;��R��MfYdX̫|_�D�B��#8���;�Vo��:n&�(:�]�xț@)�!��$wY�b�Y��
ׁ5L�o�r�Ԍ"�2����9�m+����9�OlC֋���L�ͤ�P�b� \�LɈ��q��Z��|���Qc��L���|�%׮����(�3f�L[n�B������gUL��^��f��*:��,��O<qMM�{�&a�N��?���q�"��WA{�-o`����= w��:�B�_��B�'��Oף.>V=(�
�e�Ug^���^n y�|��;�c���V�*��-����o�̙у�ܶ���Xzk� �U�m�E���
��!��f���f��%	SKx� ���ٻ����2Π��2�� ��yJ�[��@�qf��g;����n��&lͷ�g���F� �FV�ǧ♢d�VI��,	Ǫn.
H�=D��ʬ^���"�&�aL,�� =�'ж�K��Ta����}Y��Ъr�pc,Lc�}� I�`�6xֹ��)���dB%�#5P;
�?�s6�d8�Z�Ѩ��W�cK8w��D^�Z�O��h]dUD�32zg��>�Wo/���T��,a���l{�wJX�OL���e\7����߮\Y��1���<��h��_Fr�<1H��c�ǵ}������N���k��X���K�ɵ�f��oFM��߆Q�q� �&�@�ehQ�l%��F��� ��C�O�i*�[���&�'U4�-���I��'G㰟̍lH5�ʅ>u1H�����ۧ��������떳c*J�#�u\���ݬ��.VwI�mf����c�J�/�M]1�c~��+��;�8��pD�zy�K}�H�T�<h��ǀ��q���)����!�'-X�<Z�{NP	ާ�R�2��'^w�>uq�}>�T.�z�q���-�����\�q��%�uYJbs_NQ��C��t��9�)j��b��Tz�̤鳏��Uy��-�M�k����%��mb0���7��=�ab%�^��K��A���D��XA���1*��3�5�C���{ �oA�Nya4du���CώI�VN�?Y$"���a��a�^��0��M n ��ۭ��+\��Me�zCq�� ��lH�",��P�WP��?"
����.����pFԘ*E�'Hz�`� (���Թ0J��tI���[CWR�,��n�[�n�WlM�g�ί�8���$R�cu8VAdR��r7_.��
~{��@��u�w9+f���j��IQ'�
29@^��+,�RA2�+���;���t[݂�˷�F !�s�iJ���eqgk2O>b��O������iݠЃI�:� ���0/Fû��8H�O���J��A���@�a���8�v?�����w���n
A7*����q��|��q 5f��������\��+�U��fuV���^�H��'�#z���-a��A�FPB�vgn�1ӱ��@N@xC��G�W�3G��PV�=�b٩.�Q�z��p6P���6�{(}0�9T*Ɗ~[ߑ�6^�|���|���Д�u]�{����\0���O?�m(�y_�!�h.ŵ��%�CF�zN���k���o�m���Lף(�t	L�ãk]'B�U]��ZC�h$X��P�N����軂Tx��a�g�X�l]��>Q�`�9�3�V����vK�2���疓���[=���V� e�M���<��Ёk:�
#���+1��m���Z��7^�� 	+�J\ޕ �N����x"Fxvz�m������p�pbN&cO�~������sA�M�^M�>6�Ie{�X'�y�#�M"��M��䟌��/�Ƴ�dYX���Z��zY�$�4P�1�{���}�����ɢ(��W�~v�&��7��;�9<T5��S{Z��ƾ��3V��R�Bw��Z|L�<��p;�*��0Ӈ���;^�����G$�i32R=�:�̮V꼰�QĠ��S��5��a^��4�����OSk�o�x&j����҉��f'��!�N��3�Q13��@p�{��6��A���C��2�꾤;�(:������73GWC`U�0q6�A-��]|�.�,
9�6��L�6��ؔ1����R ��e�Y�.�