XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��91�����L@�*]�5͊�E�������5cK>�? 'b�L�����'a���j@�[� ��d
�.�d��e��@��̞��hO=�\�*B{b./ג�l]���&�&��������.��J������2�hP4�/���'r4�VS�`����V(�u%Vmӿ������T?��Hmd[7޷�A0����FI���c3���1cl��a& ����<B��&��ei�������WԘ4Y<t�.Hyʄ"���ʴC�`�GY@%d׽7�I��Z���ʰ�E�P���AO
$#d 9�D�}��1A�
K�j��E�UR���|x��6��u�-"��~�"���={�*�+�k>~1������R��;e-8��#�ؕ�x�*����n�q�_�1��U��±I���8���[5=8�� ��r�h�M �����>r� ���M���5� EM��<`��f��Va�h��K�;�H��&{s��)�{���Ih6��|��3��:���	�΁��/̠�J���x �~��8�)��}�]z�����(޵�NLa��?v�Ru���4���wn��UZ�3ڲ�Đk�m�hsP�����i~� qY�!a����fKb6�"��zxm�B�����r~Y���(L���84y�!)�w�f��ސ-�Rh��4�i�ɡF�ָ�&���T���|��rK� B:����/�4�A�K\=���yf�.L�l��lٵ��*1�eͻZ^��{_B�9��0%�'�bh$��XlxVHYEB    3a19     d407Ȕ�� 6u��W����u�T_��$c"����T��j=�����'�zƖ�#�����bweZ��%���!��s�p�?��%�A��Y�G�R���f�f�]T�/��z4 \�����X�\��{2��U�Ͷ(�q}*f�M�yF}�ub����x)�Ũ�n�l�Y�f��E�7@�Lf1���8��GME�珉�$��5�#]�Qgх��f)���+a��*斏�ީ��٨D��V��^���B�͛8&��e�JI��N����"B�(� ���jؓSК�e^��ͣ��yX�S�w#4|�a��#)�`y|�mm4%��A�Z?���ɀ��P����T-��
uF�(x�$��B�]�U�W��8e�Ɠ��2�_���9�Z�mH��f.�_X_�g�	�&m�nŔ��Q����~���8UF)��X%��sG��z/�Y���v1=@5X��x��u�"����rN�^��/��W|l:M ���=���w��h�r���iw�9o�t+ ��^�؀��y�A/�x$#&�ۗ��[��"�+"�&��YՕDE@��sri=�7��]��G��X6:]�[`m�Y�}��d����c�q"�lo�n�����I{�����]vP�r*[�Ƚj��Ɉ.i��)�pK(�fKצP�����A�D�-M��J�~�i�l�;΀g�dO��|����P\|���L�05��)ZL�M�Y�
.�m�i��c���x�y�Vf6�6zɹ�:�B4�މS[��5��j�.��1P��/�ڌ�8S���V���^BŮNd~9�D,�S���F��#E����X"����A��,ƙ�b��3�r�%GT�����k�$�t#Ц�݀f��҇�-R6 ��VU*%٩hњ3)�!�.�=�摽����!�q����I�e`!�3�Y(������yg(>��?��W+�����Hiծ��严�s��r�*�8��ݔ�1�H�kq�eO�f_\����l݈�Ͱ �J��,�e��r�5@#��G�1���wS2%J�@e��ln8+ c�(�1T�bT)�U�+b�*����At)H�l�!-f5LWm �׮ȍ�b1�7\dW|X}���h�`��d��M�bk�g8M����d�;4g偼ښ�W �+�H�34�;��Bky�w8� �*7tq�)+��*�_�0Y��kL��Y�%�A��7���ox��:I���Y��s�	y�b�o#���x$�)�'u��-��\��Z$'�Yq�$D��^g��7ɽ����O�>�%}�	�n�Ί��^(��|�,�ԿT>&ٵ���zG����:���
n�
^��n�WW��J�Kh� � ���aUN hI���ɸ.�u���5��QU����!��������,�(m��limTP ���q�ű��4X[�1�˘�拘����0�&��s�K��M%��;Fu�õ����s����>��'1�%H߬�w�X�7K�b��,��@=�Tr�'�h���A��!���ֈ���d���w�ǆD�ixm�A�{����3��7��V��?IV�Oώ��O_�i�0i�O��?y��#����u����L!�>�.B{7�S>͛	���@Q�ξ��_�% �\.��?>���(�E�v��)��~�ſH`�73Hi`���@�h�%Ck�/h8
�^�����n,'���o�LQ���z��T�l9|U����F� d{	�Ąc�̚d�\M���u��ˋ��N�%Ci��#:A�x��A���j�w�X���)H,�t�2n#J��ش�*�T_���(�6�:�����v�w1T�lw/[Y)�����&{V��mvçzp{���*�w��P�شKy.
'�+�N��F���B�7z�g����O5��v�U>2�_[�Ӭ��<�k����ĵ�]T"����^/�g:ӤP�Hg�T�hݕv�$k��G��$��$�ɞ×�Iٴ�H0�yx�Gq�#��}
*5��`�$��H�OV]�\Q������R�������:����U�IC<a������w��BGl!؈���&l��ŵ�{�Ld��7��������[D�����O�:��%ų�R��t�u��1o�
��+KL*���� �H��\����I����hN�%�鷭����
^ �e�����^�z��L�[XFq,�����x�:����v�w�`�lp�5N�+\����&[�ЈK���/݈of"�M����_���(e�A33?���w)�������E��;j�b���D��<��2p�m$R��<Tk|��
�hF�m�%+�/��?k�}^�^ވ+A0�����t�2Z�g��4�Q~u�[z����!�KѰ ���@���wۡ56 � !���;��6/"~5�0&C�B˛E�Qh�*j�.�K��)m��l3��+�Ѝ�o+�B�;�o�)D��Y��R���L�F�7cP�&��V�b5�%��0~��lϒ��͊T<����(J�V���[�y�U[���(���%u��t�	��M�_��̷v9*��D�hk�F��q^���A�,�$W�Bc�u!�	_c��1��a�/2 J*�|��6��-�}�:��E���^P��ыr��$]��aI�Vn�6�._���V��l�̈́Vz\5�����E3����uC��4����dV��2�l�H�=��2�u�V&a��d���o��%�?HĀ���b��
S�)��.�C�\l5�<�5����#�c) ��aP��U6�����j�2@_�aS5El<5��N�*(������K��,8����A��`���ޙW��7K_�������φ�'�@ �#ˋWt�������˻�X�m)��։!I��*���,��t3�[BZ����K���']d��])�c��*�mU>P�����No����M�T�t>�,��n �ы��W�8s�TJ�W��)��X-�L t� �L�r�s��h��аV�I��]/k�^/�XT&�o�?���Ȝ3�~���`
fU����_#;�~����k�	_s��9�A�Ҝ]!Jͻ�?bek%O��јړ��)V�"��Q����]"삲�o��5H ��v��ܧ�V�q����Cg��3T��X���S�N��bՄ7u�%��[E
"�G���j[X#����]e�d2�d���SL�u�����X����&���g�2�	�:���V���vfč�����=��tӳ_#�������r��	�cF�+��]�3��a�v(�X���N����7��b�l)��Q�]�Q���b�6F�j"�g�d��6�z��[��.���ul�5�7\}?�e=��(��J�Im��$u