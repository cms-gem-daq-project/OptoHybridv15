XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z��gVA�wV��c� 1�]��J�Π�'�e1���E��ɩ����ൾrם ���Z9�G��fo��	�5�4���4�P^C��'w������Ճ"0|yU�D�xN�۝H�zA�6(p��I<��+y��&���	��+C�*�0��p>;���Z�n�U�l�R�:��@�4Yy�Y�$Sc��a�bl:�A-&\|�9�/�&�R-�]��F��k>�E-@��p��"�x8Eԩ�1�ϻ�R.hm��#\/�g5�* \?�HA
R�?��C��H����	������e�Id�N�z�L�{n�ٷR��9R%����La?O���bN;PSU:�lҘm�B	J��	[�.^i�Z�R��!"or]8�0�e���FPw/W5�_r9��A$���`qH�+�7�Kw����E"$�`-`S;
��mYV�t��U�R�|"�A���+�3$��fLQ�^���F��x��e-�4
�m�&�v�*�U�]����`J�;r��O��� ]��EW7@�  }�ֲPN?��4�5�V~ín�$�Y?�9�!+������8��ckW�]s&0��XA��-�+��� t:�)�������c..z�b,c�1�d�ʦ	L��G2]y�_.~.z(���~����d�w�����&��ȏdZ��X��i�֝f �$���r����z�[�F٩���+Q|����,��D4�>���c�	����}6�Ѡ[��b�1�?V���R�Y��G��W�p�����Ft�a,XlxVHYEB    23f3     910΁����}G��$���[�cȹ���,���"�u��8��4Ǩ��	�3Avt9�8`n��N�������I[��#ӭ"e�Z*�K'q�<�b6��Xb�?���R0�H�Jp���kܞ�C]hY��K�Rlw��C�C\��l�$ZN���z���JI�5�̳��B�4�G��R�jcz�:7�$�Bz�Yۊ�� ��Cyb����bs�(�l+�6o��p�\���ΰ\��C\����h��E�~Q��T������|�wL�O&�""5��ri���F���f
J	�/p��1G{t�1ee4/^�E�u@�X�U��l]�y�\�ࣔ�k̿�N����C��\N��I��4����!V�e��u�:��s!�$��*�R�����p{lF�D��x@�}��u�Л(�>��z~Z<ϡ8�z�u�h�xP=i���k�q~��@w�����3�@�0#F5~��r>�X���j��.R��гO�H!��ڄ��m��%��54bb�bWۡ��7>>ա�/��	Dh
��u��ݬ��S�M�Za�H����WX�ʻl���?�D�̎�����ʪ����ŦT��Î�B�2ؼ�Z�3L�Ч�Gy!�<Q((��i�탵��ڿ�f�}��9Zb���ns�8T��5��g6-��+J��oBO�����5�,�;^'=Xx6n0���5�����J��� ��o�BB]��W���M~�a��ʍ��1�A��ՊBR���GY �M�\g����s3Qܧ�
Dx�)h�Ȱ  UU��}7Xo�R��h.'j���sTF.x=�*���R��� �\�$�8	_�|�٨+�p^RE�L��-+=|��ЧL�� ���9�9R ��(���ȑ�A��0Fo~1y�[����|Z�gabU1m�Y[��,�a+�ldeZ8<%ot&�Yy��k�33m3�R��s��ַ4LG��hF1<��-�#�w�*eKF,���Y.�!�@3#���y�á<��a�N�}�2�Wi����P���+˪�]t��v�T��X�4e�a�X�Ws�j���%��~6���a�c@3��2�)����&�T&��m�U�:�"!�[H��jTdE��m��!�Ԍ���2�P��Wo���5sI3���{���,���t%�_��"8��L�Ձ^c�ŉ�A�W����^�������p�dփ�����Kijt�݉[>'��6'��
k��Wi3v�������j���2�����5��ɦ�~��� 6K�}y�)��
}.� R%���rw�ٓw�\�c�,x�R)��q�\te*_v���A��_��}j�<�2���_����̓9�fZ�M�Ic�('�H㊚p���R��&5�r��s �R��ta��nc�������2ۍ�l^~�����]-�L���e���y2����1gO�=��S\���9�j����d0����0~5���g�+��&<�.�9\NN	�ûJNEfR9Le:vu5ASAh�׾g�	L�_��QQ��ۣ��\�(!s��me�б�-�����]�( a/����Ht+���������̡W��9Ԟ��ٔ}P8��Ej64��{d�-��Z�<)^��V~��i*rpBNװ�H��<r�?�}�x3$^��7�+` V�x���XqE�E��!ڏ\/����F'�6팱����8��`a�d!MX ����B�x=	�vDM�2��������ۘ��)����:�sB��"f˵geYR����(�	��z�JC���Ry}s�aU�v\2�=Mɒ?�E��bm��Y�Eԯ�P��z��jS\�Ӣ:Õ9�a��]~9
[/J�Hd� gr�ᝈ��4j�o�U��L����1�)M�Ѿ���f�,UJ�?oJU��=0���Φ��.�:=���(��'s��]�Z3�;n��ᐳ�_2E8�h
'~�M;.$��3d�}�F&���y��4&&��\�oB�� x=���7M��Gx}Z'��W��F��r6j���ȷX5o���x�q���:�6�N�N���k����'�T�.����㚱=��e�=���B�z/�
�/Y[�M��Q�Q�1��@a^��f����T���W@i����#g�"�#�=V8�A���r�ߠ��R��՘	O�V�/4���o�Js@m6�k��q��) "��&�ҝy�	�]�Y��%_C����|��Ȃ{���J܂,�d+& +%Q��ly�w=�|��2�\�e��R� �|���n�G1825��ѡ��&�5S����w��|���|