XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ᵔT��(����.�?3�s0�YT�E�3ｉb 	� [2e]��%��ۨ�I*�e'{�u�f�,��$px���b	�?]ą>f�.]���>cD�@Տh*i�OI����/��V��`��خ�;C��j���Y�v~hF���E���jn?<�R˹t�M6�2�n�Ĕ��IU��!",��l+��hZ�ZD�N���h;���~�}xH�&x���8�1SP���8�j�5"	��H0�g�?���VmB֩��~�"�[`����gx����]��:���j:�}FC��35��	���ok7�KdД���u&ر� #B���΃������j��"zm�ı�>�t0�#W�Q$jO�����A��ðR�NHSm�"��ÊD��M������*C~�[�X�H�DV�h��Bk�=��RO���=���k�j�?�ou�X�fEZg� �ѽ\b�]�� �yݚ>d滶�yL�p�e����P�U@�O��%5���t�F���3���.#��V�<z�h`��CwCҵ0�0������!���l�� 	�L"�5�~���GRw�X[:��Q<e2���\�ᳯ��ǯ�SH���`��݆�5Z���^���C�d3,㈬��, ��S�$d�@Yu�֖g��p��6����;���Y��He����0���9{��Lk��t��<�Q\?�1ue�Zi�`<�i�H�YL{$r����~��6�ԇ���,���w���K��b�z�������oR"#�XlxVHYEB    3a1b     d40�\	ҧi,�Ex�l�Ay7*y+/q��o�
sr
�}9~�i`�<c�aȖ��xN$��wv����<�d�>���oW^q�V�9bD罭�Ÿ|�S�����$āuȎ�x��z=e��6W/"bO�'sI�E�V/�R*۟�ń>*:�IJ��{,��\F���9�V�d����p�L���1�ꙝ���z�;(壪��G`҆���>�b��ta���9z�K�ܩ���҅@Rw;P@�J';U�E����$���������=�8dw��Ѱ�Q�\�19��qϢO��C�T���3%sN%��w	Yˉ���~�Z�k�H&�ȹ��#�b�#���V����=����Mʈ��+�2�Y�(em��]:PZ�A��V�(*$�_��O.A�n�����Kg4\V�U�J��Z�+�(�
h Ƞ�Wa���ۦ�{Cr�&V ��e��l���/$�~��NJu�EK��C>�>��h��\���0�
�h^�R]��$e��2�6;���} ��� $O'j�Z�C����N�I^�� ��a�Q�V�7>���V�TS�z�H�jU�����sb�{��W��RXM���_&��<^�[b��nJ8�6�'a�.К�w�p?%��|CZ��9��"-�T�q��EU`\+���h�,T�y�<Y�;�k�ּ��� �����CL�7��z�>�1�,��G�F2A�<�j.gGJ������+`����@h�76w�?{�3��@�՝5����2|g�*,��z�gx���ꌯ��O%G�m� 1��B���9S�e��,M��7�r�I�g�6j��H���o~~Tg��+ �/��/����p!�lJ1��(t�a��k����X���v�e�^j$\-._pv�}�S�����ˈ�gIH����P����p��j�� rJ�J�/\�ZwA㈝!z��L�����	�C#�ޚ2G�?j	�ȶ����/((�T�g�L�d>����[�Q��x�-�%��ݹ2�f�0��ؔ�� ���;t��˥a�V�@�bv?�9�]�y!q�10��d�Q0�:��})5H1&+��p �~Q�$e��5��g�kH�V2�b�b�}u��U	��nʀi��~ H-���Fכބ��~lG����)v���|R��ئ�'@$�I���iG�Å��6+>$j�7x�ʲ�|��}(�]�嘥�݃��Wu�%�h���# d��'S�L�U���c=EW�`z�� \,@�����o˫����l�V�
L�)#����J��֨����&�#{�0�S9��Cش��k��@׹K�@��O�;�L�2#�I���b���h�Н�)�l��R��%c<5���svՂ!��/)��ܛ"2�����o�"ޕ�7\�����ǋk,���.���77���麨�,����1��.
C�"k�Ï�/+@h,��ɗ#��*'����j�41�ͨ��X��G8��頩����������c����䥷Cy���5�����ʆ�t���V�*2�h̌/���0�����gS�j�˞� w���*�K���otꇔQ@@63�b>l��*�A���I?�7� �>VȘ���!�^�_�&��w2b$3�UJ�jN��Ŭ�1�I�K]�"�/|gւ�(
��P���
����r`#��r^X=Š~@a�����6�B.�9��bs���S���l�]Y\:)�m�h�a��zZ�Y��3P�䶹����τ�>]�%i���X ����	2t�Tt}к<N�Մ$\��]1��+� ��(
#jǙ�wm�rӨx����Ԯ�t���S�ZF���ta�������*rq;�~ʟ(�L�(��JH�) �{�`,��b�I�ֵjnh:��V�z�����}��;�9,]��BW����ea�@]Zp7FRQ��
��}e��c��!�zj6�(���e3&j�:����.�M�[�`�e����S-�X�G�lY��K0��H2�<���y
�� X2��Q��F����ˏ먜��CK6<>&�`��su]B��q���!`�6��+��$�AJ���:��YP�-�W`
��o^M�h�"&��2&�>*�d��@G�0�"3���}>=�"�;�������߯))wt�-R���I��D�}0_9��|��!F�����ٰN���8M�w��+�t��fH#��jG�}�k���	���Ǌ�}]ղ�簢B�Y�Lƶ���B�Η?D;��c-x1��[��7�|�=���]�~��<
��uJ2��}�3��C �̶5���(�����kDy�*8�.)�#)	�7\[�,�Kw�����B�Ci?��0��#�]�oj���z���4�6�n� �%�+�b	G�LNR�8�Q��3�6*���r2�ӢEPD^�%Pc �l�|�
K� VJ1��y@4~fcݠ=���wnլ����5��ĳ��Hu|�j��� ׳Q�S(b�n���eЌ��F!���LY|��?���H���.��	23��.H-,M�Z`�b���T���C�Q6X5��F�!��~��bR�匌NwJ�$fb�ʿ���g]]�G̮���$Ty��+]��/�s�&n{*����(N@���3��r��9<d�Þ���2�����e������P�
/��SM��.��=�|��qI�����f�P��a�6���:4���LO�=��4%�ǥ��r��ވY���G��g�����P�H��gڤ�kI�j��
�=��K@����[G��Ռ�jG�~:�W����KD��#��͓_���7IR�H�)�<
�P�=x�Հ��������EAu1~�>h�g�K��b{^O��$L�Z��̇�6�D
����K�he)��tCb2L�${�TCN@�qGpmKu��%��ݓ�B���ɿFCʮ4v��)��bf^k���LAH�ZB��z��ދIn�1�L�Bs�M�ӌ9uF3��(���֒؟��[X���
� �(��ՍY��!ŝ�E��5m���<�cK����$r��!hB$���0��j9�ѥ���k )[=X�R�U��w>Ts�����mn���Cp3�R��*=�^���|Z�S�N~�}�CA�<���XE+R �
� v�E�LǬ�[��z����\~��r�_'3u�!K��!/vJ�d3�O���B��=���=���h���w;7/�h�d�D��#m�=�&�e�\ᤂ����f$E�<ל<��M�{�2�\ (!���f�p��qN*�%���q!y��o�|"���5���iM��z?���^�(���FHR�@�0�,�)#�.͚��[E�_K��&�[��z�gV���"gf@�