XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?��kU�N�څ����!�*w�=��ک���ݻ!���`r(�Ɠx�aF�
r���P���DV��˪���"���>�w��v>+��]�����+�H� ɂ�.B�_{����m(3dx7���cxfu��2����:q�?$!u���-{v~�L&:N�:����h0��-������Gn�6���������p�U�Y0l��_?�$JX����VIwu�Д�E�W� ^r�N_�u�׈��C�,�6�����s&@� �Ne�������n8�����<���!rZ#���E���AG��0��wO��0�w��!c�Q�u��w,�wH��u�+(�SBaDp�>q��M�R�ǿ������U��9���ڳ��m���y���qk aι�:wɠ�Kg_���5Lፘ�ꚽ6E{|�"q��E9�u�+=X�HXo�����#�!D�La8e���Ƙ�=Д��S�}��vŇ���?�:$v��-�������b���K�7m`''c����$l�_�o<ʻ����향��@px6�H����h_s��D�@��+�[�t�;�h�ɭFz�K=Ib��'���K 0��&�6���ʥ��UF^A���	����vOd+��W#,�.ߣ�#��I��r�4'�ˤ���1꙳�T�a����\�Ze�#e���Xf�d��C�u?�����dy3n�����ّLA��^@)��Ǣ4��+�m5�8�l�s�ǡ���V~�<��yXlxVHYEB    41b6     c40">劻U��eY/Ҭ���Ia�I`��z_o¾!�	�߄���7�,�H������ �
�,�z�#�=�5b�4^ߊ�ʻ��VB��k��o3o�F��Q4����΁u^�E4RŲ��?= H%�k�D�]=}l���na������׳�H��|�o�0���k4�}Z2��W�W��\3r,��^�s��9�����4n>�9�:f��m��!�UI��/��y�U�jH�"#�'��وXQ�ð
������N��P��d�6WO1DS��@1PO�$iR4 
���r#��7X�ڭ,�^Y�e��$-<kA��&�JYm�������A�����E�&�5�s)+OXg�Ȧ6jP��@�'�s��\
�O'�T?y,ZU�˙���+&f,�񄸖����Y�����F��eӛ�'��VK�AQb��E�4�Є�����qd�ֺ�I}cǵH��бJ&�YL�n;���z��ɿ��08(#��HO����Ⱥ&N����+�&�|�J�_JX�e�R)��x��/?�٬��
@�"�H5��9��)f��)�c�\߉�C�wg���)���a�-��1Ӕ���8YW���܄GVtYS���X�h��j�=3l��ŀ��,eV8VS�Me��l�x��X�l��ۨ9��3 �5�jw)�N�(���@��-��d�U���WU�C��R�?Do�v������\��X�npY��h�Ƃ�ZAM5�`���Y�1��x9�pQ��⦹`�01�o��ß֫�eUɘw����c0��2��Q�Px�Xbd�R'(z�s@�*�$�D�T(h˕�|��!�"�����UJ�ށE�c*m�ՠ�n����Wv	�b"��������t�?��~u�>D��S'J�������q- �o-�[��u~q�q�#D�`��f���[��}�/��Z�=
�2�͙��'�^$ʗH)[-��W��qb��Bܭ�G�ʡ�?n�TB�Q���.::�Z��	8OUz�GHۿ��`:s���$A�8���C_Q
Y?b����`%Jd�L�M#��S���g�xW9�&s@��Y�a5b����cc���p_#��&]&�N`�qR�Ǳ�j�4��d�����ű��`��97�W�g��PG?-�c��@��%� �Aa��	lS���):��?�2"H�/���CBϸ���C���8��F��o66pA�G�
��V�"�O~�S����1����h�z5�ǵ�L�z[��que��%�ry�_s�P� ���N���#�eQ5�΄鹌Q�	6�t4�x����¼��0��W�ku^���)�UkyԹ������J��B�yD���d�8�Իo�gpx
����w������IW�"r��p꘣�W���j�!���%3�����ˊ�����+!���]&8Xk�nY��5�Gv"k���YH#ȋ��+|�u,λAt�7��)+Aq���#�S�D
Ž�S%p�|v��~���z���U��}C�7����u" ��]����zFh�������H�E�Z*��(v�%��P,;0���Y朝
�C-<�D�:�)�,���|��G�f���wJ"܌�L���_��3���z"���G��K�E[�
%�Mw��'j�	3;E,d���k����ZE��I��t�7b5;�V�ۺ��a�� �b��]D�	C�Ek?���(�?&Gx�d�Ι��! �0PRW�'x$ uّP��ˁ;p��\7=o�о�)��g�G��6�(�Z+0kB������W��� ����}	�^ǜ���v�2�X�5�.�X���-��*d�T��d�p.���&	�Rz����8��{#T���{YN q�]���r6���V��l��[x�+e ��6�&�}1���I}���6�N�� ��EV�>�5T�I>k?��c�
C�#(�Y���p� ���Īw�:">�Z2��p��	p"Dͼf�_�	��� ��*tl�ںi�8؆�m8�qے�C�v��DB�Q��F�NsT�7f���}}�N�jp�c����1��=�R���=hk��;�_����w����V1�X��h^���;E��C���S0�nQL]��I�3�u����~��,�����t���[�&�����G���ĝ l �������f���ӭw�Z)��i�J�UG�?��?�������)}T���ɜ z�����C��Qހl��N���Z�����C�Ouѡ`��z#��B 2�(���0w_�6r%�h�����?o�2�x���BW���O��&�D(��")���/�@��ls'��B�}�MU98�wk��^��1�!;?/�8��'�r�M��J�T�h����n�B* �8��YH�i����e��?r�����Ӭx3l�G<�����$Q1�^�{�("�����K���&���p��T�j^�f�։V�b���|�(�?E�n�}�$����k-zݜW�|Nɫ�~�M�91
����1[�JTY���H����5�X��R!md���/�hM:�B[9����,�e��.O�ъ����wq�B��>����Q��w�b�㐮A~e�v���џ�J�,�->;������(˭W�`�$�YS)��P�|�S�׋>6Z���*C�}^���<W��S���MƳ�o��4��*s���G�c۳5�tjg����̺\� s����UR��p�53�)?�Ȋq�j�gv��!'�,����P�gz���W�X%79��.1�z.=� q�?|t&KG
UJ9�Ln$H�f߁�+��e<���]yT�-�8�D�-�T_/3E'��ԃ�,�p��Wvf�p1�-�KJcb�S��=/�u�ŭ�x����PE��S��V��A�xݫ �r%��n�V7j��.�@���|��{�㸙r�TgS[��թ�+���;��:~�f+*Զd{f+�$�U�u
x	Q��/�hLS��@�f�X(�i"�`�cä�|S�ޅ�j�g��݉ly$e���~H]������C/����~}�-���1��⣅�U76%8�QFw�