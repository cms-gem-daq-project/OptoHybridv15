XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����~$�M�`N d(���m��o-R$�ش��B����Âne���*.�[]�H�ك�)>}]���E�`����Y�c��$]w�����N��F�����-x�լ��ی� �Fh�?��7T�\�FhH���d6�H��ްA��*k:m�x;0�(S�]���oÞʙ���Ow�
�����N�Ტ�^����'���϶�i�Q2۸�w�K��DA�do����)���S*j��&r�XQi|��R�+���Jn��^[�U��ʦ�fQ�*{*z�Fw�x��6:%�#��G니T}AQ�6O���5�L]���{ȕ����������&<��֦�Ch�ňi�˹��gƇ�՚�l�rvϖ�3I՗ΰ�Ht��F��	�����e���N����rúuە1���1�h��Ĺݏ_�b��}�
�6����S�s��~�\}yDp��!r�s�R�f�߱!6��5�s1�wV�'2�7�G.(��d�~�+�E&�Q�ʝ$Y����ɗI!>���j� ��ݸ���ꍖ�N쁙*���1�(l�7x,m�5�� �C9�� )���ysI�M�G��ʑ�qfz�WA�����	��d�#��OB���*���j��� �@qk�+������t����憀5&�O�=2��=HQ����6��ݺ5��s����p� v��ɪj:4��	2�C��$��/�F�s�D���������^%�o�? G��	�*Z˲w����H�u��ʔuOa)����F�k�uS���i�XlxVHYEB    4e25     d70Z��x15k�x���Bũ��8S/`�����Fn���2ʝ>ޚ"^����o�c�)�����8�3\u�M׭����@����=��J����v�L��hJ���*]��G�Zj��U(ɲ����u� ڐC/{��]Php� �Pf�n��/���(,��{�$t�/��>�,���1(�vef����n�����k�����4z�b;��w����	���H�x����`-�զ�\���Az?y�$pQPwٮ��㤊"pn/rriv�K���}ui0����1��\E���ozb��#)�>�߈I`�3�ןB�;&��S
���
U�:����ۈ�5�n���]M�u/9T�¦g̭E#)V��A�z���@p\�C���6���^$=J���Mp�)K/8�����n���o�����'���Z;��9^���r���5u^@aÇW�ի��
b�-bI�����7!�2C�a���A�ܒ8'�	��X�y;C�׎�g��oI�~gD��Ս���v[��$6�H`�F��h�и���`#�F	:�e7�Z@��ł�q�%���lt�Y�����Xݧ���G.�
���/ԇW�Ȏ)Y�hw��;���~eT}���73|w��J�)�����m R�,���%�%�0�N�/Uc3h�m�>�p�JyPIj�O��G�#�O���'NWvF���[w�,��K �ܖ.��؃����~�1 l�8U�Ab������n�&��ST�7z8F7\*�Oʌj���EI��ң�ǉ��C�F��z�����[�C>@�nDb�K	_W�K<٧UQ1�V�xv�ii��~�E���#�ei)a�ED0����7���B��7bԖ���s���`�P	�F��Ny;I�%�S�٤عpF1�+7Q�E�v$�}U4|Z��yl����=�M�+TvZ�״"J6�F5����T���[�_���ؤ�o,7}��)�$����;���Z��xs
��z=F4������H,p�^f�ß��@�ߓ���7�^�]��h|P�<�^%�!c�	���X��2��;Ĳ+�+�T����|4D�4�7��ReX7ۢ+��A�F��`�G'�i����p��a��ͤ�j�qJ��#��|���C|;�����(U7�x�V9y`�u�f @`�G(��LJ h?�|[�i��<k�kc8�� �#U�4t,a�����)�!yzc��[&����`���V[^(�&34��!LJJ'mc(�L����N9ͯݻ���Q���Vإ�]�J� ���R��8y��O�iŒ�kG�U9?��A�?*��ʣx+�ڍ7�Ib9@G9����`�,+��~̤w�RB��Ï�4ø��"9�a�W���q����}�+N31g������%��e�G9�3�,<�Asc
��a�nr�׀,_<����=P:���w�W�{�lC��,�bnتU�Ғ����(ux5?�f-�X`v� �7��N������j4��X)z�=g�����������0& ����)�(Nr����u�#��5�݉_�ZW�S�Dn�H�c��rR>���W�»�D���n�3O`��P{ҸRq7�����`viӑ��v�� ��M�}�|1����Ry��^ʇ�B$.���ڮ1a��<�9b�%���F����'M�Y�3�4~k�/y�P��oU��s�s_L����6<�%gh.�k�a������-��ih:zu��v�vE�RR.����z����
�5����&���x��%;���:�����t~9�9͂;���!-
���?�K|�Jc2��^O��B� iSV�C��gŹ���������G�����=�]A�X�����QD��$������8.#���7�����7�7��R)��r�+�[��Bv��v�(�I����@j��9iAO��f��`C$Ѕ�����=َ޼\�A����ՁM����h��Tr�Ċ��=aY9�
���&V�<��K=����P�0� vk�q@�峱b����ݛx^D���L�j���ix���Q��Ǥژs4��sx��9�ǘ?���]Y'�l���n=$��~H�V�� 5��e��,�.F��F�ɫ�]g�� Л��_@�z؋F`7���8����Q���j8}S�Q�A#JY�p1�d����]�[��/���'tր�Ai�-�^co�up�US��]��܉aq�aN��]�����י�,|���������Wz̑&�'Іi8gNL��~,R�dҭ����;|1=��"�gE�ƃ
�zph%��)e�W�Fu��=P��I��?�Mȫ��k��t��J��vf��}�?������6��� {�јr�0Fa<>�n%��n�>~�3��i��Ze�F�Y�b�f~�����?�2�bz�QX�ĥ譢�+j-�<�f�H�x��,-��z�}
:ŧ��q�>��5b�p�J+t�񋸺GLn�&�h����p8q��ުԷ�oV3��<V/Fq���޷4����M��	�}��X��$����N$V	7B�� }61����Φ�����`:�Fz�'N�D�����rN����ˮ��a�~��fzƂ�4-�ש���ʂy�
zi�X��O�2d���	�!�!���ߛ��C�wLQ����X�Q�zլ��ȉW3�� .Ǥ�Z|�,���M�����_�y���[2.ݞ(�ڦ�T���J�.�ĸ�p�%su�Oh<�1��bV��8\�0wT�"�}�a&8�႐��!�qȆ_�'U�nD.Ҩ5��Uգ�߇Uh�Y�Q�Xq�/�@>G�a̠槂 �S���	�v�?c�U�8�
�l�D9�q����;��k��Ȏ$����%��//�@�B�G��P�[W�-1�Q	������AÅN�*Mp�N����y�i����Ї�%V}�8��ՠ���Gb'�u�$&�?�
(S����/ryqQz���a���Һ�Ń�8�i��E�FX����Z�v��0oJ�Q(%N?op�o�9��Ó4�8�'�������R��^'͋��������o߱flV�~k<+������ߣѽ���g�_���p�^.;[�Ȇn	��fO��_h՚��ݍ��N�~p�NR������������C 17μP��w�;��m�Pi}M�r�~b+�M��F�Ђ<F����?���u�ކ�ܺ2�n�G#NN�{�*��� D�uf�)�� +x�P�������'��=3j2cXN�0%H=0{��s�%�P��`Σ	ؤ��\��3�,��kW6��ePܐ�p��<T�r��^TFXw1_T{�V���&���t?N�	�՛�J)<>�w,��B?rܳC�u}B�Ո��f�����R��4츻�j�U��RzL��g�