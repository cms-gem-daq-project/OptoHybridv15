XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J���7���in��`���B�B�����cd�tc��}�=�ގH��N�"،.71�hs��d���J����*�6�� ���E��=��jC1y?)��xI�}�B�%�V拳͗I>�l���Ȭ[���%g�H��=v�&̈́��$L�P�܋��t���Ρ�#�Eم�6�:l��A	��I���K�v��PUw�C(��.ͤ��#��B�w��'�|P����8"Y����8�]/9��+I���F�` 67+rW�	�{HOq�ߊ���*KH��c�I�C.��;����H t��+�u�t���^�}���pB8P@����LD����6L�S��&{� �8՝�&_�{�VO΢�D�(���˩���Z\e�W����SwuZR�Y�M�L�Y�4�Č���a'��5�E�H�{U]4����~�ule���2rSI|m҆���/7)���/k��6�
�1�L�D��.�@w��"3{�!�LL�J�@��m�Yl��FE���f��yQbђ�w�D �d��t�  �9�Ⱦ��o�([� P�ϣ��7���l)�3!���\�0p~�~2�`�H���d���o��	5?�7A�o�,����I D�/�7��ҴAv�ι&��RLv?����VPB�R��{	�B]7���h���dO�#�S.�mwS�&�T���M���&Ǩݵ�)�3����vt����[-"�u��Ĕ89ް��l�0Lq�w7E'ܗpf�( Kk�}XlxVHYEB     9e2     330����,��pm��n�;�:��ܑw�#���i���S2s"���LC��D���B+`�Q��Č��{O&�a�,�Q�c�&�MN�]�"�D�UO�$A�{O~.�X��J#�SQp�R��ۨ(�埋�6����&&�	�_�B��>����9�� ��\aP���l�`���Ϳ�ʠ�V�,8FZ���=Ù��`#�ԣ ���LT��[I�Y.�;�#�D�ٮs�ߡi�b\;���V��P9DpX.m�p�U.=�<��<a�R'�K^��܃��Q�����~�T�R��3埸�>U�`�#-f�Hn���5��KԚ;���Xvl#��s�C\��.�vwg����y=j�AH����/��@g�#�F���%�#x�|���.v�+=�?2>�ևjơ���؋ ��g&4�T�"����CWXK�|�R\ݢ���&�D��2?���?Akv��>������)��-U�]PÏ<>� �2�G�>�m8����,�:g��Xi����8���+����!eLzo6u"/8R���@s�!��d���)Q3;:��"��z� ."��".9�R�����Dnb�i���M�҃ۥx��6��-��}0�M�h1����b����K�I���<��y;�H��a��jd��#E��f5�ض%�4�Ȩa�}4��CO���F�:�B�>��[�@�9=��� �(�����D�y1Ԓ����7��:D~2ʧv0�6�����zFU�C��$�O7�]WY��H]�J;:�@��3���F�ܳƹg���D��ƘJRv� h�