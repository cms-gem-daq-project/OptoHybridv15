XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��yk�[2�*B�2�ڨ-
7K�JD�<��Xs!�� ���Fh-<W��.FH�
�����<,x��SBV�"�{�JT����Z�R���>O�JUN��۹
��T��=�iifR�vw �^>�Ϲ���[we!Dc6�MGB��9$:��'e����L� ������;���3���$�NNJ�Y�3,�B��m޵:�M���M+��O���m��l��?��}� ^�/�d���0��=	������O?��r�� ��-�����r]�#L��C�l=�,F�7G�&���RH\夕�X��9\-� �鱝}�"��#b����.�!)"��RȇFL+������Q�8�����m� �.e�?ֱӃ@J@������"�����Tަ�M�IX`x`�N�'��R���n[;����3�M��-i��,�BeC$����{weƑyL}e}����4
�r�F�nB!�WBpl��Uvo5Ӫ�#�MD���/��Eȶ��y��T��5��2��/���%��K�F�kO�1ưr9�k�-��_!���16�o�HL��<�4��ѳ&�Z�G�9Zq�������.II7�8*��A�Y*a>7����Wv��aWU-t(R�qӳ�NE�������"Z��D�=�������R��6������ВU}D�[�m\����t`nO�9 ��m}��Κ7�S�[
u-q7$#���ɢ��a%�~�Ŗ��]grB:��4��U<0��^�KyVC��/�>XlxVHYEB    3c92     900'�aH�2��^h����7rXOon��y=j�r����V
eV��u�!���I򐭌�@j~�с���iF��if��`֘�?M�Z��� sj2���a<<����"�ϑ��~>ϫa�i8]$ȚC�?�����.-@5 �b+���*�IĔ7	iT�����]�oQv��1��h��]
R���Id��fކ���>H��������`����_��98E"Z�ky�{��0�p�"��z���GXviֶ��Nq$w�9)�ZȎΖ����yQ�q�ىn��1}�Ն_��H�iܰ����i��X��
R7LBO�u��3C�d����Jh6���=��(�O�E���oŉ(+WZp� nV��1����)�Pe��>�!�+��e�|pX�����U�<�l߳�5'�i����k֥�~G5����pua�J�y�#����0�R?�6�\�iő�:Dv�[9ۯ���W�I����ߟ�"k�|	@�
�j;�5%�=�-~�M^�@���2��-E�}�8�F��6�W�=UEl�=���=�G�I�V{F���q
0�jU?�h�Re��-���;�H�)JBL��ҫ���
�����O4��d[���;�}�w��0A�"Lj��O�c�DnDU4�Z'��%!1��;]	jD�ݝ.�PX%4DR�R\�e�"Au֯l�W=	gH��<�� ��'��?�8T=��+�����n�P4����%��a�gR�12BM�+�|�Ѹ5B!,}�t�c��_v��g��&�󗮔L5� ���r�+����ϊS8���� h���P�z0�A�ޙ ���JS�����À:-o XrxGKո&����� Ϯ�9�F;m�xb����42���+}:��Zc���;1��r����c(*ܷ;L(fB�������͛��:	n��l	���V�ޗ�z����no:^�i�L��(�l�_�����A8|N<�~�4&X������OSc���,�"��5����|
�8,Z(�q}x����v��q�UEca"� t'Йx܆��/��� <�;����[" Uw�ɭ=��[����`�i�~]��L=��|"d�;'=��O����*�SI�P3�7�=7 W�a/�i���"G������m\>*��C,��:�ϱVo
�s�M�h�,�؃D7�}�⍋�<�h)֩lI�l�Qv	<-��F��yV}�D��[m��.նB}�Q��]:͍r�^B����q�������%�Kq�s���$B�L�E]�s�a�m��o�q{�J�h�p/m^q։��U�B�I#�dMLʴ�����:m����T�yy��/�*��R퐓�-� ����.0��#�\���Q,ț�hW���,����z:�y����-��7�˼xfdzՄ�	玱�N�9e3��R��T`X���1�����ĜrKO��k��Z؅֍'�����e�1�DIG^n�N��7����:�6�	
o�����o���(М/���v���IW~��S�{�z}5�Ղ~T!@���w�0����A��t��@S�R���|U�Ƞ.����;�=�!35�;V�YuS�N�s��tI������~f��cƁSО iCHy�U��,�Ŋ~8K��AO�V��y:R�����,}�o���P���T��n[2��o�ˣ@*��0*�0�i�X"�2/@6>t������F��m�5P��/�־h�����[*�q�U��kW��#�.�4�S���2êe�{9�#���;�~H{�.싯0t%<��|���v�����W��O�ᾥ��_:@_�b�/n�GkV2�NIԓe�*ᬁ�M���
J�>�:�;�B\دq�6|�w��q"Ht@E�(Z���"z��f�
`�[��b�T�u5U����(�i�U�����4,���丰O��<���?8��KՓ��P�wb�dF�����R�Z���=#R��D����=\g3V��l]�#��KV�z�7��Ӏlg���+�2�{��ǒ

5�����M5^c�ys�����}�ѓ �9������B�s���q���_�*���P��ʡ+�����0�r2a�|?J���K��>��v9Ѻ6�[1�#�MW����˘A��3t�=�E[˰,=H߰c��� �\PSi��Ui�'��:�',��}�K��4�V��^�Oԅk�~�!�Mm��=p�@���#�R.�ԅ�X$䙮R߄ƶ��Pъq_���*�.8r蟢�A��vQ]X��u�b����������	p�<U�