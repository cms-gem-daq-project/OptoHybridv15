XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��4J��TWw���b��x�nߑX��F��T������V�"j O����3� _����R5�Q%m�hs���h���FfN#��EYo���(C�$�+����Ḝ:2F�-���D���a(Of�I$�N8tt�u�׿���2�F�"�]� fK�9�ۡA��`L�G��$r7�S
浻,�b���U¹kW�B�r^'[��z����^@��u��q;itW��Е�y�7j�jgh6yVR6�:Qb{�gl8J6��;����΁8zE�B���q�o2<U��O�$ۚ�8����gz���b�<�j�6�lŢ�j�Ybs�(M^_wF��ON��;����G��Az�t0�T��u�[� ���*\������1%Zp{��ի@�|�C���^�00[�P 1L���瑈WX���x�u�c�5����d�ǂ�A����|9�2u P�z����[L��nW6��)�}�����3��m,����2�g��z����Fӝ,O3���̥]|�ĔEr�{���8;��T^�G���2��� <����x���8�x2A(�S���\;�w3���'�<N�q>��$Q�s���R��Ζ�$�9S��jJԥ��g����\WNfmZ�,���u_�`�5�h�$��~pR�2 tA,ͺ3z�����m��Bv�v�:�a&:3��s��H�-����K�U:2ڏ������f���L���U,�(���U��qW̜NWXlxVHYEB    38f0     d30���:p�hm�Z��Eq_���L���K,��B�?��@���;,<��p�@a���h��?�ǠĆ��u��֕L�@I�=��ʦ�����8�N3$���=�?��rq��<��*<PAv�#{���Wf]���86v�3���Q�L,��(�䮀�ꨠ���Z�Uе!La�����Y9��U|�)����D#B~M~��ɽ ��!�<�ȗ_��U�l����kɃ���Y�lqᒀ�\��&�I���Cv����:����&B�Pfg�0�R]|N�a[�ń����Vkݰ깸i6�y��Bf�1a�R�R��1�1�$΅�H��8ē������[9(j�v�����־�H�,ݐyl�_G&�F�8��j�BΫt��H����3�ʶ�%V*�p+���	'�[-k��S�~U�#�v, �+.t"���S����>gO�[�ŕ��[���j����Oz������i�K8Uє�����
�Y9�;c���b�>��{)�l����'49$xrV9(�Y��i.^����Fv�F��F�V��@Չ�P���C���t���02���0_��D��ɺmn� |an�����R�{>�ʟN�%�h9���+�`����G���vi��}���0Į+�����N��rH
�ю���9k9���o��=��M���@Z ���%	TCbNs�2���_�Y|^�J�^*8s��X���ݓ�	#S�KO%�$ww	��w�Rl�0r���O�#�yJ��;�\���yӘ����ZIi������yN�Ja����]�搢�P�I�sa
�TFN
u�V-� ���;E�&�|Z���2�s	�����B.�h�_/�-���m�@W������"�)J6�Mt�I�.�pb�b�ϳ�	�ޟ�Zۧ*2�η��M(1��&v?[�0h��\D�s=r%��O�J��W��Hlh>�]�W gp���?%h~3�%��~�87�d�8$7�5g`�Sڎ���J�/����>y��^���e�-��ɾ�FW�!��4�sy\	�Q⌓���_�/ m�8f72쾓�\��(.x]�R��`q���C��R����.�U�|qa�Fd�qD����[5N�wDX��RQ����o�K�Y�\7����Yi�+�L�)֙he��X|D{��MP]�s�4Dܞ�xjr�d��������:B�~o>�zz�f?����)�)�H�J$�
�x �{���BS�/ �����sK8�Y�y�d��?�K8��5��8,8i{9*D�P��)�tj�4>k�4��%�]~^r˩�BT�~k��vt:WvW��u	� #���/P���d�s<�!��ޑ�g�.�]����z�'���� ���$��lHb�� �`o��F���w��,�8gŌ�Dx1w�f�?��nKs���a����͘vN^�I�o���tlD���7/�Ӟ�L.�b�g�����X�-��8�<+�X)g~OKz�H���l���"�
�F�׬E���
:�Z���*����Q7­2��[�(jE1� ̗��P�g$��>�a��Zt�Ц�H�t�#�Lvo�����gnm��!��Yz�9��ۼrY���D�Df���R�������(����U9}�̖Kf:=�Q��%	�׊�Q�@m�X��@�UA�-J��Ƽ�襤~A]�&��@���vJ�<3���Q�)�)y��ҿ����G�\��w�1�������߸v�>�^�FoIx�:
�������#�E���!㱎�|�G {3a��b�0�Qf�\^R�vH ��������_�?}��*2��VaC��ho�}A,<�}/��� �(����;pX�xC^ʌr#>�j��3u��5�E�|g����G�gH*(�.9n���K����g� e�n�v�O#R�.�W��&�����I�d4�)w
�i�7m ru1m��XS$?%v��U� k%��x�9Sc����_�o����П�(V�z����V��B�g�㽧I�ˎVJLDq�.q��p�'���/ ���n8��L�|:Ka]!�% �c]S<˽��4�"�SD��M8�h!$�^I�����S0�}����
��#~dc�����ia<T��OW~i��Z��F��ݥ�v{�i[���� x�S���Y��t��.b`(�1Y�c>N)�[ڷ.uT�;C}���$�!�lCN�, ~[�
�eKeSl����?D��Љ1��J|�vrش���{�]ɸӧk-�N�!��mE1�:�%%�!\*e0�C/���U��,dq�z&��l��*%�5���z�z~����l��c���6DR�F��{1�BȜnau����&��/OЮ2<�����`D[�GN:����ƇK%�T@Y�[�ѲhTBt&u}ez2��L�7��� }cN���.�_�H�b^I��^�����푓���(�3u��8�T�b��D��GWuKs�v�o<,�ɻJ S�3�+EKe�)�Sx�U�%N�����l+��l��~����<�R! �2$��o%CzrAg�=���k���i�=���e�U�iX˴�6�cЏ�=On1�5���p���n�Xuo��`_nMm��d�?0�����a^q�Zm�:��C#�v�h���+��i�M`.���b�й�[�pq�8�M1j�'���S6w)�\Z�}�I��͸��=Ў�Vf)���f���C�lƆ��<��V�.~�2z47�������v�,�_�:�i��M���/L��M�R,�܇��"q��/��0*�ݓm�M�2=�.:��Q�6F?|N֌)O�ć��y5-V���I?g[tV�eYo9�Ww������$�Ň� �a{y�Ӻ���-�8*OХ�/l���i
��k3�@������1XCKǣ�nD�ir ����H�	/�ת67�4�7:�����fE��|��(p�y����)}q������=)cZA ��]�p29�$q�}��h b��	/FZur���>1\'%2�=��������j�����u��
�+*j�k�~��bG��<q�>O���[���|*�v,g��X��d�
���ĝ�Hm����#x�ܷw�-���꧰_��1,iv�*7��W"X�ϸn���C���h����CpB���Z+��O����0��Ҝ����*���Z�"�W�����w�}~	La���ɚ�üo�g��j�K*��7���_��a�52u" �]��8��?��%E�Ix,�-��.k	���8�X��b
}�z#P�y�Rcs�G��G������X�>2��B�?+�j	�}˃��L��'c��Ҭ5�}�E�\=�>�$�����H��������TQ�'Ÿ$E �k-w��i^���g����)u�