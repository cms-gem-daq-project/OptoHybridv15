XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����n�SezL��O>�M/��o�v3�R]��G�k�]�0f�����%�<��OD`�s��]����t˅?��|�L��LDqA1�d���e�pk�לu���hUy(2��������<�@��|Wg�$jy;Ok��IҒ���"ɥ`&��mi:�ܗ�c-�9�F3�@���XHfWt��R(�e�<�,1�ٲ���%U�bN�߫����ȥR#��~YA�	�F����d�w��(���2�l�d��u��V���*��Y��AmlO�&�}L�џ���N����.n��g\ڡuy*���'_|�8��	?H�C��X���W0�x�J�9�ꛓt����ܽY�o�����=t���II:0����VV�	����YL~�$�SRݰ�>&��.���n"�����D��)Ӹд�G�C���`���r�(�/ׄ�쾧���y���{��oo���ܶM�Ut0׊,�=s����6������+��jn1��'�����F���W|��z-y&����pF�61��Q ����f1�z���0n�hnޙ�G�Lt�����{�5aPL!�e��/�����E�Z�N��ZPWR���c�����Į���K�a�_��hJ�&|�M���ϥ��$x>�~\�� ��Z�e��+pa5B~sM{��=`tF��9t-�}���X�c/�cIf'�餕o4A*�Be��-�8��I���q�:=����`߉�q ��c�3S'NY�erxB\���j�������A.�U�Y�_�XlxVHYEB     99f     360�؄�z�D�4�I�>;��$����KB}�ң��#��<����E9ʅ2�X��h��C`�a����;A��sK�����o�<͢��b�mO�8��Mo����-����+}s0�9r��d�R�5K,���wňy��܉^Q|��<���!���v?�G��ˎ�i35XP�����ǚ{Aǥ�4���+��e�w{D�>�"���c��r�H����Mp�P?����拍&
�YXS�_��m���㘦m�I�G�JO�QС�6^�$��a���	|_"ZvHfw�͊���և��(=lI��P��OEht�~��4���,tt��l^��ɑs���ZD9��Xx�ebj������	,��p!T���j#����2l����L���`W�@�{η(V�f���k����ǝ���%����Ë�b��%�2��}D�X������`�O���uq�O��{\(pF��+O&�L�x���;H~����).gFxCr�g�!ѥ��t��0W�#���TV��K�-t���^皉'��j�cG�6ԙ��,�<�����c"�3�D��>�XW�@��|�o�X2�s��j&:�5]����?�m�{���!�] r�+b�X��GP�����>��̈g��u'�m�%�c��G��9����@�K	�ET��AxRG����E��nRΏ��)SR�2_V�?0>��8��ϣ�S�w>R ݶ��d:Go����1��y-d������Q������
߀LlÕ�>����eޝ�kFG���@$ߩ@H��A�^�A�x� ��'��D�Lg{X�V�B�����}vO"<gD!��Q���n6j����5�