XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� Θ�����C԰�:����`ς�a��\�
�
�s�*����J�[��4��Ǫ��x���|����6��*~Q0Sw�i$�w	Mx��vmgp�CEr����CJ�@m@��u�&��x3hp3BW�΃���\��|X��`���޹��`����c$�@��Q#����۶|�Q��l��ǔ���*m^�̓0��֤��/�n�{1�b�_C�ٵ;���
�ȟ�q���x�U*N5i��*#I�h�^���mrҎ��ƒGuN<}{��||����
vo�'}�Ѥ+#�ʧ���p ��l�x�R֠�d�z ?�W��	�]4-�uV���CJDoR'	v�b��29�-E�.�4������C��EWXf����Er���D����]�4�@����[�Y7��l-�(�P�I���&ڶL4�=	��%�v���"���$��d��8�=j�����ۢ����G	���=��C����5�d��M�o�+A4>�
Vk�V��@�%��N�+ϵKO�/V�I��T^/�g�E���+%�:�w�y�Pf<C3���ޛ@�G�$ZYn�,G���@O�2D�%�2*�K�.{�A%E �B����������hN5�`��Ֆ���{;��;P��.Cտ �4�2��߳dfTd���`d��K��D������nL}�Ǜ� ��ŋ���LJO�v��W�|�@Č�����B�v{�C�T£��&���_W�Z�Q�E�I�ϳ�*x-�~��c8�x�XlxVHYEB    d88b    1610IܡZ,ڔ���'Og��ΰ�Q��a�@ه$���l��t�':X|eX "��!�� �c+�ڻ��׆�%�#����[G��&�zy��#8�Cc�'d[�"^�Ch �tحyӲ���aE�C�N�`k	�W�fpkpG��
Q�B)��4��O��_0�_���O	��,|+-�]e3����2?zQeO�-UJ��:�/y^e$iB��5�*p"7ʊ!^�;+�"t�y':�  �[����m�u�{�������U��CP�M��oy)͟�B�P\���� �@c�z\���HJkYbVdMgk���V\27�\�J|,�o;��,ı����-�~H���4R�+�R���Wk� kmX��J����5�(�]��Ľ&�ɹ��Gwi�t���1�hk��[�p��(rQ���偭��k�:�a������`GU�,��t���ov�Z��@g��&�mfHa�\��h9�I77�xp^�������Gr��T�q{�6�"��^�E+���b7�)�Af���K|��ݕ[e�:(���[�;t�ǥ(�$`]S�`����	���{e 8�)kma��VR���/�$d!͐難�v!1�E4��ǩ�F�q�z�g�j|~E\����Ò6��Fт jq�aDYm=J�mg�F��lC�:����8���4ܱw�f�ľ\�
���q�B���#}!��+��NQ����%YNpt5<����S�`������%��j�Y��+���&�g>��� �1}��9{P2eMF����re}��ޙb���KΣ��[g���֝b�E;���(�]K�r�t��h�G4ү��A[)�莔�[�:�n7O�k�X
3�`��=Mk�6?�i�%�y�ƹc� ��h:����Xy���n���A7î=?F)
���v�CwN���6���S��� ���� ��t�i�K�H�z�5gۏ�2p���P�t�&�?��J���J��Ɏ�,�j���`-��)�4��=/2��߰1V�9v����zV�[�g�x� ��=g�Z��t�4E�O}���aX)�=��2���cc�Q���7݁V�����ʙ����WK��b�o���f��u�֔��
�m�a�0��2=O<�C��*T���8��a��wߏ5� ��g�g%�� }��R;�gC�Q�O��pM�F2����(ͱ>f�i�Y����C݃.�H��U�6Z4�k�NX��֗��2����UP��9������l}��i��k�-*��A�	�V˫wY�Mi��~c�0��h�sԱ����)�%�����`��:�?N�1�MB��4�\���`ʗ�0����xR��VGN잋O0n#��#>��e�G|2G�:�d�^��Zʱ,�k,��`߾��3���[&��>�P� ����M�`�&[c���a7-y
�O��˳T_��-x�➥����P*x�.41� ֵ��wU"B�w=��~e/x�)�F��)^�-ĵ ,��J ������	�(���_��^��6y�R=�jݣ�@����-����v�p��ac�*�tXp�w��?~�ˮ
n ���SX����K$M�"���)��� �cq�z�f��¸�
�W���ga�㚂?S��e�^'g�˗�H3@uw�Q�q_:�A��L@<�r];��ʓ���%������,����l7>�P��S����aۋ�_>I⛧�ֻy�P�b?[ЋH'<~�3�f��^[���eP����Ũ���H�+�õӬ���	��M�M:9o;�~&_�:���t-�o�y�4-|�/:��%)4È�v���9G�
�@1�J2Gn�m�,m<�U e�,6� )5�u��[EӞ@�Tu	�h�Xx�1�K)�T�w�?�I���0�G������l2�{��"91��soE��}����Һd�P6�@"p��1��cK3��l��]V'/G|"��(��)��1-Y@��T���w���k��؇X�c8r�k�c�*�EN"�<�bng�T(��H�6�+�-Q��jɗ ��jǮ�޺u�@����b���؈�ׅ >�M�G➯��^�k/co���	�µ����Q%P5�p&�O4�K�g%��hi��3�1#@D�:���3&=�e��!K��?,ϧ7�R�j���|�]rS`��[�`A��S�>
��Y���w��`r��<ؓ�u�G ��b��/&43"𛺸./����T[��_�a�_�Oj�+I�vS${x���U���[�z�$ye֏�ʡ��a�ULI��:p������y7���ɒ�1������h�>�_)і$��|=�\�u�5U�C{�ޔ�4?"�����q  ���hLӢB>p_�Y;�)�7��Za\>��fJ7�h5��բ�f�?5�'A��u}.i�Y�)�Oᎇ*�IC��U�\�[i���zj�#zJǿv
�rSQ�f�۱xT'\S��@�4�~�]1LuR�g�)�__�PV�E����\=sK�h1\�k݁;v�s�>3�u�M�s!�D��D�q�1)��E ȇ�B���/^:�4��B�b��H\�t[m.؉E:!/3�7y��Px��͜ӱ�DA����&�Z���%��<�7�B�f3v1�}�FB����Z���̀�_�f{S� G�S���fЂ�|,_��l^��A��k���H�Ek�[%Y��[y�P�6�+0��LZ�X�2��v���+@c#:�~ ��~�N[Ӵ�V`Eв��A���G���R:W���#���_�.�.G�'mg�N��#�u�4f���$|P�����i������3B���a��s%E�H�'PMJ�w���弔����B�����x-ǘ0���Ο8vj{��;��og��r,j��`(���Ҟ:^ȫ���>%=ׅ�|x�]wA�I���m73����<�`��,D�"��&l:lF8����S�чҲ8���	��^N���}��CET����3�vp���:�H gE�L��$_`�E��&�m�]#T	�)4wV�z3�ϙ�F�+��W^r�n��������}yt��D:���:�i� 5W=����6I�6���3�_������-���vN&��)��i�{R��|c��ڽ��|Ο�d����'����P3@�'U�L
!oN��	Ϲ`k[��7���[aW ��e�:�bl*���6���;�Z}L�7;L
|oe�b���s�����ʇC�6��)w�s���z<cpQ#ްp����2|)\?X @ϡq�A8�f�Q����Axe���*/��W�~~I	�	�l���pi��+�h-x�{'�����6,ʃ#�?���*��0+�挥�Һ���Yod�s/���B<+�أxqs�,�8LC����3A�w*¶[��2o��d �6�X@+��{�)[dc���� ����CR@��T��&�f �bF��9�~����u,�P:|���U^�����R��E� �:��f�|��R'�[wn�^���V�P��7��<b+�L�-VIN�	�-��*�Ϳ�߁d�,�TO)�"䱷�N��=F��>���Xr�'�?�fo��L�Ef5��"�β �>�[�l�)�^��%}�!�U��.ז��ӹ�P�VtU��i�򖕰��A��e�{Ď�+E��J�t���j�J���N��|B��9]���z;2-ȽI�{�9nڃ��fM1GP� ��6�
�����z�n��jG�7�W�CƋe� ����L�Df���h= �_��o���+~:U��5�!I��̼�0S��!'��&)Ur{���s^�2�<�]�	�N޳�8��@C0��Y]��l7�Mp�x?�M�h���v�@�xB��-c��3�b�ۚÇ��˰7�9�\�1�I�Mο�n�<s�|D�������ˏ�)X�,ZM���x��$�日a�	�:���1i0����\3"�>\2�
p&]֮��b�ț�K� ���Y�����^�rT"MC3�7B��T`����'j�I��8��w`ղ���p'V,����WX��x�SH}�,� ����@Ąr��8��߯���L? ^�Vƻf�c:$,�A`���o%��f���ɡ�cιx�����i��cl�|Bqg�{!�6��':��?������ `���=˚n�#K�O���'!���O�P����H�;tPۜ�o��_\�4~#>��=����4�;ї=h�R���هao��G�=C�ȶ������#�7�: ��3\犡sX�R|�Mi�9�J�\1��uAhyu�m��]��+��K�F���:��L�5mЛ��e�2��v{n)Q~�!M�Y��`��K��!�'�#�������%�Ј�\�@��©�p�Z`,��J+݂�Q�S�e�h3l�*Ƈ�e��D`��֘� ���]��,PL�3���k(m�>��u�f��ݮ>�Q��)Y?'�R-��o�����Ǒk(Z� �T�)�A�#h�%��V�3��*�{�Ҿ��8{��3Y�@ ����;�垤`湃��Rӝ�˃��0�`�K��J��<���+�P#p�@�4�%+��G���IT���a�N١��:��
�ƽ- �w�EkT���'b�" QHĭ�����V��o7�,]����?��b��&H��<.����+��>�b~�kY�C������e�2�0Dfp�~x|4������^ʗ���e:DZ�)PH�%���fIw�����S���%���zY��O��T��[9`�O��E���ಈ��-�����Z�	Og!<ƕB�oT�������Q���Y��wi��E�λkU��2��@��8�oPk~�E��^F����;-�c���7��؇��{�T��EK9���nc�yOc���l󻐠�kM�iѬ�!��J�&��I��neچ�.z���_ʤ�����Wp��2�td=��	Gf �oy��r-�T!C��
x7��*YW�Rҹ��W��UJ�;����yϙ%�3�5	�"Hv[�����8k�^PG�v�\ŋ&��A,��,j��ď\gE&��}��rpZ(���L�Ӌ�-����#��	{.����r�	�Z&�D������9�`�z�����R�a�;D��PL�r�$�I�	;��xys�7&�C#���F<��7���Ҡ��po�,�	Ff�sXL�~02zU�#L)�����0�څ��v��x�H�g�B���N�O�*5� `��@���%V�j�3���N�$�Qc���7*ڧ�p���N�8?���H�!�U�DJt��(u�W8��x�A�ot�������M9�|y�? �b�M���uw�������t2�5f�F�H��ݸ���2 &ZΥ	üM��I��-֡�8�-.��E����oRq\�ϲ	��S�!M֔TF��I�GG��H�bw��T]Ci/8�>���Ñ�����lP�_c�
�t��us-~��=�!ɜ��o)��A�mb�E(�\�r�}E�!eTl�h��^�����D�����>��DͰ;#"0Y�eY����*\x�Xo��+��8huњ������6��Yֽ� r��V�?����W��5�)�kWB