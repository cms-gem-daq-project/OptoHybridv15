XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����	�@���D�=��i�=V��VUaZ�{.�<���;����'�<���o�<�	K�ժ�����s�5@K����|M�����
MW���I�y¥�]
��D��P�ߦ�Z6�������Q(�rkn���V<.M�����9�(�<.ѕR�n�]��wx8Л�$�6�cњ�]�bEU�	
�8%;��x�	���!M:�{�5V��'�g��B�5�����m�]�U�̣pC�'tc0�C2�{$�8�-�[-���=J7���Ĕ嵧��H���_ϣ����u[��tb;�E��O��+�[m�-��8�#�/~Q����w�n�0~m�N�1��	U8߿��{=~W�J��T[���<�%.�Z�ʣI��M=I�y6��Vv��&���8c����5�l��P{c�t��6wړ�'��c�K���qN±�`؂r�Ac�܇���ނ[$�lD9C�[5��j���Jz�Q��!�v��$�'�Q�0���	��x�ۏ���8
�?��s��&��y�׿J^e�Ú{�ȸ��E�V���������'5��c��d�U��L�Ma&�pp�������j2��.z$2�e�� 6]����~f�LM*<���x����HI�����GkH9�7��>'�9���Ru �.H����/�<�P�	���-`��о�	Ox����u��:�}4b������VN����*_�C��uE�����VU#�@GwpL�H^~�x������d�j6%�-�&M؅|��t
XlxVHYEB    edab    1ad0sdE�����h�S�_��FU#z�SM�X��|K ��s�0��n�Qd�4l*&�-�W�=�Һ-	�}�<P��'6R�2I~	��;�/�7lh�>�ɿ��K|�n�oH��0�XJ~���Y�E{A xׅG{)]��a��$��A��b���3�x����L�a��w�j�����%0�`tƎ	�o.$�ҳX��I����%�C�㜖&0�p���c�kxfH�5��k���\L��BӪ�����C��I�5t ;m�Z'G� ��'�D�^*����SW���/jx4b�u�����e�a!���+͎��W��R���;-
�?O��=�AP<T�5K�u��.�J���h�mavXr���9�hh;�$,hh�^���@d�\�c���|�[�5Ƚ��/5Zh���{A����P��s���m�;�� N����ksl4��t�ܖ�b����c���[���"Y���7'�+�dͦ܎�b����n�2V�%�]p(e��b���qӕM'�w<L�'�2��'ץ�@�I}�L'����x����5/tp���,�I��v�c�+���MGtKTu�k�zj�e3�nC~�nh��C/P!b��z�0.�ͻ!j�{M�O��������HO;����&_=ڿ�>&r3:6�	 ��M1�o`G���k�6��1g3C�o9.���7�N�"bl��rfE�=04$�������M��z%gX�fFu�^�S�ULc�r}\"�ރ �S=~PIJ2rxoGdً�Un�����/=��#t\]����%���(nܕ�Lj9����ئ&��~hЮ$h�~�J���i�>���U��]\� �[X&4�L�G��5����P% ^���(��suxsd��$����\���QB�W>��3�]d)�F��	Ie��p�7>DT4❪ӆ+���D�˽f��
�����÷,p&w��B��gLM�����a$pCQz�yf}2-��1d�r�7��m�ɖR:���Ȋ��1 ��~*@rԇ���9���O�PE꜕���O;�A*Ӽ�f�DL��̣��􅷓��K�wX�e��P�����]L�:._���� ��wL��?��&��X��N!��U=�l��SZ�:�@��Z~YS6CSlN���֥�u�|`W�n��c�[�s���������]\�E`�$��,ǋU�����ߛ�	��n����}�����ԏ�^���BQ�d[	 NlA��Fu�����ܓj�@�[`I ��||��W7�T?��-je���ei/��W����Vl�ޯT����m�I��HGF� �p�C[��S$��$�YC�_I��)��޷���S�Y����{���EL*�h��&VC�����A/�kg���|��p��r�A���}���M��`�Gk\��42�L�����Ӂv�o���i�,�������9%!!�}
5��C�ل���	���-6��ϴ��<!��G'&�?�_>2b (;��Tr=��M�K��	p�T~�?o�#���
Ǌ�w��Y��T�Ҙdu&7lGb,^s'|p�/��3	�����h<1u�-�ݲ��VA��!\���c�h���1����@|͜pن4�n П�Q�y��A�qt�����FӬөW�\�Y�����i���`xIϫ�V�i�{!�Xq�!M�E�\�rr�[`���I��9An{�M�XCЫ~�2^��T}ާljR�yZla0Su�酺,#���7F�¡�K��O�||�p�����Ѕ�b{��lqP�� +��H���w��
����+�͵�l�K�ֳ�N\���*���ջ<�s܄�B��A���Uְ�#͔�C�z'�a#��Rb��pE�R���xy^��7G\y�8�q9Z�bL��@Cސe��/�-��m�L͛q�v���p`��o��bbk`PH���ml5��w�����u��dF�]*��#:�s�u�KIJ$���ShY����|���v�k�C-�Q�d �zy��y��٩BB�42�@��oE����6b}ͅ ��%��4.����[�JT����SǕ�-J��P���[�m��%�*�NPW�QX�[Ы�ȩ�c=mU'���O���""�R.�#Ts�vѰ�Φ�PXER���|τ�����������um�[`�Ǘ�d<T莉���E������$�'9��2�0)�m�k��u-�
�k��'��Og�e��|B2]
�|���������(��b;4�B5�(�k��~30Af�Ꟍ�	&1�ڰ�?��}K��l<^���,�D�����\�5\nǠ��b0s_�t�f��d��e#�o^v�-��*�ǥC��9;��#��:����9�jB+Q�����!��E��u�D^9��j 5����fS�I��B_ߠsA^xGZR%ڴ�V=I�?5U�(�*�w��։���vT�'^�]�y�����ɬ�b��G���^~�9��a�*n�w�����L�85���9��3����d�K��ا�p�T�0��*�hfQ%)
��=Ii�(a��ojq�	u:�O�4��&�a!BWJ T��K��i�qy�L�O�_�d`���
�.��L�G�)�쨿��TcW�׻j8��
��f$t �=KoT{̀��▶��8�_���Z���\�e�x��'����J���D��'��v�ܲr!�~j���ںR�.Ͷ>��2�R*��<pN�(��S�W� /� AM6�6Ѕ�J����Z}�Rv����	���o��}7�� &!�>�'a�Ʃ}��"b���&��E�ѣF�6D��T%K[���[�K��,�o���P.J a�j?�����G�I�{�&�FW]{�X�ĵ�ۯ��j��E���t-����#�	؝�sx4��c�Ϗi���q�F�z�~����3b2�����+Vxŵ�#V����������yt��r����5�N�h�Sy ǻ��<���C��V����T	�nA.ÙnhߝZ��/�E��������?�h?[޵5M|E&ny<�θ���z)�����*�b��Ύ%f���`Ur�7����Q���`��j��bIi����<�S�\�V�W@��U	�L�c�Z]��co�=1<��c�#ZI�'XP���[bwFuۡ!��ѫ�D�@�
pyU���c�����#k�݌Y4��<
J�*��d�y�*�3�-*�zD_��ˍ�J]kw�1l�����l ��伫P�rhx����\�e�a;�?ݫX0�s�$� ;�Le��>3���F��� ����'�{́�qb	ZQ��f��ǎaoay�����}|�ME/�� ���WZ-�LAIJx�$2�`CIG��y5�@!���$Ϛݡ9�.��9��v4\��j�&��Q7U��_ʯ�).���@�.���+/-���3�(C�3^��p�LBݎ��Yw�Ne��L�%~�Qr��m=rv�?h��_S*ڕ6��VwTa<��չSB��`/&�
wu^�e�__�-�cf�T�Q#������F��X�f���6W���zß��N�k	a+��h��ّ?|�B�鿢UX��_��_�]�&�11'�Z�;��
"��f�f�SZ��"���U0����~��[wG�b']������	+�gF�҉n��xϿ}�4����K����G^����� aZ���C��eQ���m�D3��&0v07���x�����E>��;U	)��[�s���qG����nR��,�=���ev,��wcC�
f��I�_+�c��5���1Й�L�@2�>4��UB�8뤨��feG([Q�q�i�XϢ�>Z�l�z��R�&/�j�U?�&�B0)�L�����su��Yh��e�k<F=��q�Q�1[Ã�#pS�!S&��1zQNwVܒ�V��Ǫi��8��5���>�O��������d-"O�,�v�4���~��d6�%
:!��W9!�������β�=�R��U��uw5u�`��=�&�X�����Y}�^��S6ㆰ�nJ�����=������=�f��k�ڂ9��F}kJk�샃�ۺ�g��_�#�I�=�(I�9�����t���*��p�5�Y��O�i�bB���@o���q�y(���±�ݒ�\!pqX�pڬ9Ӕ�E
�)!M<@��]�/t�j *���79!8��D�JCYo�hvj�$%�ҩ��<ˋ	PA|�Ԋ�<#]�6�N�i����#�&gd�>3��'���� �}B���ާ�%�����p~f�Ee���j�]:�#��kT������5���]�t
ˆ��~�2=�PH��N*��q�c[~E����BR��ͩ�bȀYz�Nw���`A�g��K�@�vLI����a>x������
�jmR��*�=���٫�0]�֚���o1|���xn�'�>@�#�8/�>Sl�L߲w�`BSۯ8��D�ϸ;%RCM~q���~��q]���^��^NM�mɿc��!j*$W��;�A��+h
.���BZ���[�� �u��I�[�ks-̴���A F�k��A��b�K����	��S !$�n6�3:i��ń��'����|[��7����51}��%�f<�p�x��ΜώY�HO�-p�/��&��$n�EC�d�̡�m�
J�S��7�_-���3�r�1�Q�#��#�`�}�''�K��>�Vi7��[3����Ħ
����d!7��g��/�Xc�(}��R�g֊�$b$ԿX����2��_BTpt�g%��g�\��X���W����T����W�GϬ�ǹx�����%e7s�����)]��}�f��ڊ���t�EA@�a�� �_��C%�J�D�^3)�j^�]�1���&'R9��1����M%(�].2yD���Z��P��:��t��'Y�����΍P�^�BI��
�}�b�q>��^rsp��% w�k��-���L�eTu���.H�{k_ML^����W��1�*��E����TB�:d����f�<�3��E��t]C�8��LP��pz)�X�/����!�f�T���M�?�+�sL�G�d4l:����kH@((~�{�x )�#��&l)3=8�Mn�{����f�^�;����g��3�-ٮxNf��ؠ:�E���W��d�O<]��O�������	-�|8�2��R����u�{핾RD<����{"��]#�)JYs���Hj��g�/2� 7��U1���rv�k^ŀ�/�ߍ�s���Nz�-p�V��*�F���eP���=i��{*@�p�Uڬ"L�y�(?��N�"A�60#��LK���ph�.G���SZ`�w�~Cݍ�\@�&lngl�O&�� ŘzcCh !�@(�z�o��j�f^�cv(;�Y��$pQ��za�D�J�-*�����s���+���x�����-�r�hQK;�2�0
����x�qq;�ǃ�N�;a�o;�bц;�{fD��w����W�j�9Lᘆ>�7)һ��j�g�yO��rE�y.� �P9 zF�ܵ���m�� .��fS���j��0��He[[�\<2�$@���Q���\L��xoUj�����j��*b��Y����~�搦�P�@.�U��J�iS�;��1��Fj~�a��jJnJ4�Y5�2����zW�٭������Y�L`�x��	� &<�H}�{G3}v��TٙH{΃�jn�ro��$��h�'�������Qx��:�x?<iki�9�sM��/�o��b�i��������˺�����-G���d
"f(�I�IF��C����Y5�K7��xML��~�yJEk8���(��~;9R�J��~�&�0��W���J��CD���� ͸�e+Aa�k�/��x��x�s��?,�򺼑�����T�_|�g`�P=�����G��1)�n�����zTP�HAg�s��sϙ���H���<���~�<h
 鳕�Go��o�a����/P��,E��L�V����-I������v�ӪE}�s�=�`��~�H˻,�Jͷb��m{�����-�2c��]��8���ܜ�F�b����	��܌�yԧ���`c>h�,��?H�k��Y�."�)��lCۖ�%R㜭�È]�aI�:č¦��,��_>�]vp����ѫ82���c)W�"��%!-�BpzE�S�3䌶��qm�Cɡ$ �9f��K��a�lQ�1EpT��4�i����$ߔ� ��:3ǂ���+wzdS1�-�{��k�v�A�����t��"c?������)C�*�(��x������|��P��e�T�6��V9��6�h��#�	;�t.���Mu"�F��Y��k��!���D{A&��5��Ҳ<>�������_&E��J[�W��D�"���DW�5�,\��=1��d瀍�*���7���H�}`�6�+:��wu�������ߌD���7f4���q!mV���NR?+`�궕��4���D�+���� ����X�8����yfLk�_|؃��{�Ĕ��~.��s+y�(�)Â1q�'�d]�g�\,c��~= ���3Y��P�F�^T��������}*�������rI� 1���YN�~�7�f����C��	ay,t�|PI�GZ�+�;o�	I�����FK`����"�E*����>t	�.	��nc���h��&-��]�ƙ@[9!����ȑ