XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]��YS�yH��Y�����ѡ?t.�����غ�Vg�)���7qȈK`;k�᤟J�~^��7���<n��9�A���S���+��0
JB?>������z��pÇ����P�Ux�,-���c}�U�\��=v|����.n�����'�ּ?���V��!��la�01�b�P4(�]r�g����H���-�W��sC{d�~��5�_a/w�E$���5M�?:��VM�y�5'樬��������l/R_z�GnWA�0��͗���au�G�a��X�Tt�E��Be�:�ٚö�p$8��R#�U�&�)$?Բo� ������!���v�3QA���E�B!�fx���p}82&{L{���J���j���{�lt!wE� ���SǥJO�=�/R48��`��>�¤Ty�������G�]h�U1����=� ���`�����F,��I���[��%baȎ�&��>�s!�hI&�N�=���$ab>��weoZ�K�oi)t�yr�u��*�}JYy���2 >و����1$��#��z��p��ʉ�EC=�F��͘�f2<�(p����<�g���w�������@�[|o S`te׌��	���Ⱦ����{@�A�,�˧<��9p#c��Y��)��8YX9�ĵ]x�1��G��F&t�5�R1q�垇T`��.qU�N�r�?���Zp��(�z��A���D��r�����L�t�3��5���X�F�^7R�K��XlxVHYEB    1047     4a0��涞�
���V�S����
�@��mXd�%�lh��V���f�?�5��(���Z=�=�''�Fn�>q��,?k{����]�I��h��Cۮ�%�)�&�rn����!g�Q��A�.�q���lY�l�05�"��L�����ʚ�_�2$aΑ����l��Ăz��
֘&Y���V���-(4���B�3	k0�Ƥ�M���iQX�Wҽ^��\��_��_�@���G�7r������'��7�6H=M%�@*�ek�c�Dq�'��ޢ1mt�hB�8�O~8�;-�s�x�x��=5Q����j�NH,|�,�d�	-5xQ�v=*U�^^�^�8�M$}�_sJm�f�+7.�|k|��]��Qb��	)���={��k	Q/f�;n4)yc4�ޒ�)ݧ���+��)�ɘ��x4,��D�0�0}֛�?"~���Yr�9(]4��G�*���l���Y[��pKI�<��W��A��^bo����k|�<(�KY���Ei�~XdQ�7�o�M���;C�!��2��Z�:�.� �
MJF�,a����W�\�4.�'����
�V���&ҝ�o�݃I&�,����T򻺔�:sҵ[�܂6:2j_>Hp�N�)灄#��d��bA��m�?[��� oM��5���\�>o湯�ެ�& ��Nk�	��[�ч��R,J���z3�8S ��1�Q��/�N_����烬y���(�K)�]d��{���c�w~6-�-��,��[����Q��UB4���H��b�4�f|�r���D����^7_��˦7�����ݲ�\ȃl�������P���9�\�D�H-\��D�r�r�2�#W��*����S_���T�ʦ.V�z�#�~��^t8�<]�%�Q��Hn4�J��@�z��[��3Ųj�c
���0_�~�Xs��̺�$�C.�a��C��9\*x\O�׷�y����ۣ�`u�3U�B��XJ���j��"���O ��MR��"P�s�[������J��^�M��w���F���^Y'M������;x.�p��q ���IK�3W跒�P]�S>�Vq�D�5��650��d��\��[�<�l���KoHI�2Q�{���+%Y��w��[�����Ŀu��7R=�ӯ���Ƀk�i�[;��