XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D�i{Π~�(�!���|����d:4w��~�r۞�=���� �e�b�� G�$a�`��o���`��d�l_h/�ђN�V���-s(y�^��[fXT�t��_1�(�+��{�u<}�t�,���s̢x\�#%?�����ܨX������#�[{g��%j4�:�A�� �A?�W̐!5�����i�O1�K��_����T�d��K�0�8�����Th6��2�c8$���Ŷ�T�D3{�G~���PD����g�{�4�t���`Y����'6��`�$�CB
��2_�q�Fay�2Q>�y��'��MYbA��W�A߷Rh��X��P#EcƩAK�B����o@#x@�wiK+>����n��y �����)9���~���d�������� -�|M���0@�r����@R� p�F@�'��x<�z���F���W��e֜x��g�Y`���S�L�8�wՔ\)�t�>�c��HPwlN�	&�ɣוּ��j'oB�M����?�fZ��ߝ�8Y�	�}Iٵ����"`~Ա4xA�����j�'��J�=!�Ȍ[͛#�|���P����3�z/�_��V�f�ˤ��p�D���6�4���+��?�~�Q^���Hq�ז��}war�6�<�,��r��|��/d.�z�}�r<�VjV�E�r��cb�Ka���/��39F'�0 ��m]q�w���N:����i��B[�k��ߜ��*������ *Y;��;���b�k�����N�
qhM��XlxVHYEB     6c5     3006�`L��-�9��M�)A> Xu�XaY2;�S|A;�e�ZS�'�"i�����B��#��ˈ��g,�������Y> hl���
�4u����ґ��0ȹ�r#����B$��@)�n�
�����M@��օ!���@��a�(S�����Q���������pyXMR�+����tl��N��}������D��;�gg����؀95�[�Xt��h���$�n�ܸ ��ȵ�D<�|�pv+����F�:�S8I�YX����m,p[�m����Ss��W�� :�:ǭ�%R5*��ٸ������>�����R]%�@PL�"��"�0��!���5,�@�Ԑy�-Q�c�e7J�F�����:�|�mRBQ�N�����6Pڿ��P"�۲�l��8&� ��.�5��	�|��5���;�m;��
�0f~�E��~*Re�$�����"�hy�B�HK��4�F-瀤 �cL�Nڇ�.��<��/gpZ�[n+��g��O�*��˲�ѡ�W���x����yſ���czM��H2�Æ�48;�pR�#�W6F3V�]������-�P������:��������E���Tn�t���.\��f��r���ٝ0s���'"0�5H��9<u����?v�7�+�����J@HS�����������yXK�����aqDB �/4Ag:r�5G_�I���Bq�j�
Mo����w�:�� ��C���
�8 m�)�ͬ�M