XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l��]�c��B�;e˵�t\� �����
m=8����PA'i9���B�����A�;�'ޠ҂m�n\A�A&6a��q��=�_����Ԗ|�6C[D�'�`Y�= ��ۢl�`�`C<U}��
��Ĵ����M!�Uƀv���Ə����n�3Hz�G�p�EG�����лy�:�Q7�ay�[_�p�Ldٺ�IN�O)Ok�n��GzMF��w�_���e6�z�Y?΋�1}A�#�����	�� �K�Դ��C�~��ώ9�L�| ����¯�h18�B���q U"�����W�t'��`���;���_b��rMa�ZKw �J���Z��C��Wh`�t��z�ys:-�Ã�E_��_
c�茶�?shW�@���~���D�s�T}���x3���$D`�t, ��؟�C��H���G�&��)�?[	��fk-O�����v�}�Sτ��:�&N������=M!����~�)R�s(@��Wۙ
��/��?�)@,�n3�#�����d'�o�]���չ����`�q���`�%g�o��n09B���֝��=��	��:"ʝ� Ö�B�]�ĚMI)�lHvOׄˉ���P�X��	�����<��W��t���aTa�s�X1ٸ����!i^X��Z|?Юr����ӤSO���qB͓(.�����`. pP`�I2`:�[��N	���ZYw3&N��!׼���L���":�	4n��v!�Z:u�1��n#������x��զm.a:�w�XlxVHYEB    10f5     490N�-���I!���@p��`ಱ���� ��!R"��[�?
���[�4����༸�˭�kiS�h)�möZx����.� �����������Բ����>y����;� �m
H�eZIwD,홗%�Ԟg~�ޢYc/Ŷ9܁��(���z=�A,_U��o\R�k����!�L�sn����:+�&�YE�qh�+��R��qq��=X�]�2�A�۴�%�;�����xA��	.�zc�K�F��,Z��<[c��q��t�,V�a���a��*���0o���f�X�?%�pNU�_0�7h{�+ɷxˬ��s�%[�j	�
��4�~��0U�q�z���V%&��K|~-p�.\I:����6{�m����2�aw�f��W���ZD��n�oH�<��[����Ժ��âO�9�;��߹e�Յ�Fv'��Se2BҦ #���_QE��ʭ~�nrh�ո?Xj{��jT��[ݲ��x�A�����b��}.�X�7�d��v����nY��D�M� M�����T�/�`��y߯-����.�
���ez|�n$� Hd�j��Ppw�ܿ�f�u�X�Ǩ����R\\X٩�KA(��ȄI�GX�<ο'�WN<N��y���	��"��2��ίH�S�b'J�{"rD�V �����^:8+pvX�����v��4�ꐉ��X´��SHSq�����i�����0�Zka	�@����������op���l��[5�o�P�3��z${����T|ɧ�Ȭ�1ɤ`�5���u�.��ֱB���L��3�����u�4�1���9}�$oD(JU/ʞ��w��R�:�F<t�3�j�3џ�5��������)|�I�C���xf/��O=&���4
\����)�u2e�Xnp��=�J�jʪ"�b&	&����P"�p|�F�/�r�i�_X��F5���>6^�|Nsa���B�5�?uʃ	%#�����0m�&��" 
I�/��N�*}-0��2wP_�=d��4ϛ��=*u��~Cc��T7F���2�ƙ��]̢��![��X��`1!+�
��l��?�5��z�0�sG�x��Pw�����<!bX�F�hw�$��K�0*�f_\�7�
�K�mD{�t�u0g=NbL[̓�/�~+���@7���{t>@O�h��u~��y