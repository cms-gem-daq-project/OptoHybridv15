XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�Y��^�%���Cz�
/��ί��x���iA�
�DP��o�%K獠��aD�o�����h���}Y��s��A~��g��g��+���Wb'+��W1#J��"w�����I%��7�u�u���=D7��U�����Ŗe(��!�ۜ�D���R8�C�nҫ;��e���٢�<㤍e��[5"7w�t02.���L�ac´Xc [�����33�ξd����!f!V���!H�JLQ��m�R1����c�ݼ���N������ԋ����J���aĔ�3�QB����u�� �
��?;n.r��̎lr˒��x��Զ�Q0�Q4�q��H�Q���7-��7��{�lT����0'��Z���<��k�����yH�'�w�;���}�#U�_�� >��u�|�Wp��s��1_Rh��(/*N؂����?Xp4[���Q��ѣQ�!.��n]%��s��_0cd-Z�l���%�fN���)%h���O�ԡL���x/>�z4moƣ��2��`�$ܚ����Š�,j��Q�5W��k%$�Ay�̝0��xš(Q�D�v�8�y��ܛVlB�&��pjt|����F�rA��ZG<��xv�L��fd}��]��ӷ"<�`LJ,�w�&d���7��V�8�h��O-�@��!�롳ɭ?�S[F�����F6.��@�Sөn��Q�fz3���i�ۨ����$~�7�z��q��|s\��tYN�B�����=�Pº%XlxVHYEB     7d5     300Yb��%�/WE��06y�~J0ټ��"�|�v��tR�tr��)��N�D6�d�${���k,=��v����Y�>ğ��UHbБ��9t��\lܓ�.4�Uʊ��Yx���*Q�,��އ�:���NI�B۪'�����U�`��&V8��W2(�O�����Jf�:���g|b�~a�gne�ex�<I$�����Wh�GK(x�_���	ۿ��+�"'��_\΀���+�l���!`��r?�2z���<����7\��r5�N����Q��W���4r�_n͛�9��x�����w��Ȝ�F������O�[p��x�#h	�\sϰ��jX	W情c\/�=Ǫ��9l��f�ew*���C=���=K���*V����#�;ڦb���Fu��LB��WE����OO����|'^��IV�;W#������^J�a�:�)?&��d����L��O�hC�rb��Q?�#��'3�����;�<ʨ��ldc��gXN(oL��/mƕ���ޮ����Џ��Cv�g�T��m���z��}� @V���Ѵm�&I����21���	����n�
yr1ka\�y�:if"u�L���X�]ƞ� @ŭ�9DxF��G��;�R��q�/k�����Zo3� �
rb+�]
*P_�'��z��'��젻�Md@b�u�o,b5-��Q\Р�fF5�y?�ow��i�ls�N¿��+3��b��4~ʷ�)�d�Ax<ؗ���滭�$#����S��m