XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,R*M��״�"��wnsh�~�3�@�'��a��q�!�n��ѕ�Yϝ_Q������ ūҤ� ٹ?T� ~�q,�7	�������:_��m�ˏ�.f��w0����u�h,+\N�T;��I5�UPA�!�:x<�sz-��HN*&���tt�c�}��zR�P��CU������p�@ [(���/K��rH契�@b�mW�6�y�JY?
��K/u[)�ZA����X�?)�2�"(�qތ��!�GT߭�Ǣ}=�}
�?��棜H�b�7����>���q��Q����Dhb���,ac��*�$c�ŝ� H4�b����|��*�1�=��ۇr�^��,�髋k��|�������A�`�)����7���ڮB�{����`���9ɒ�I�����d����\����
Mz<=#$�H���>0F�[y��Ȝ��3��I�D
&~��2;����aa��������I1��S�������es�?gJ�"Г,�/�m8���������ё�i�+Al������_#f@Qښ�#+��M�~2��+Z��@$v��@ZT�8%�q�×��7'ۀ�c����=a�v�̗ �B� ��[�����PM�Z��-0�ْ�_�m@q���/�M\=���km�[o,�8�|T;l��6;��q����o�V��/��r=x�<��X�W�B�L�n���\���u1E�p�th�hO���U�_5�� 6�"it��^�qF�s�Bv�1w���w�XlxVHYEB    1569     590���z(N�Is:�E�����L�"U�y�¿�ӱ�da�>����U��M�^���TP��zӅS��Βo�Gx*6�W���r�@XO^/�"�h�*�O	AB�l���!�.�m�ex�(��rS��7����K$H.�XCb|�����L^/ls���me�΂fC8˞-ięI+����g���`8>-�3�������W�ǡy9L�s]1����
�<���{.���P��cL�x��j~;q�L�`sZ�B�T�
��
�K1�K���*�K�M����'�}��r�&��ǩ y^��Ae�-�C���WL8�W��^�]�#�O�'=����{ 2;�9��bvB8$+������Cz]�!0}/���P�`V
��AE�ƪǩ<=�~H(ϧ�}�	��t@rNs��iG.����~�!ܻ��_�����ϼI}��!s�)q�y6NuVJ��%����LV��5�5��L�;��E��r��~Z�R���X0����չ{� �9���r��Q;eW�6JW�ɶ�ؘ�$a6T�X�x��%
���\*��߶�C�����B:�h�F�����Z�1���]�l�1EXy�#U��Z����>�0�|t�Ѡ�6�{H���k�,���������7?�e�L�*��T앛�`�a�|��U�<X���d!��i`P���"�L�+�����qb��Lȣs���_�І���
�~�LwlsQSR�`J4��H�N//��:���];�X���S^r��]ת��<��2rL9FM0�6ӷ0�V��PThk
V��O������{k�*,����j���֥WÛ�xq�q�:����4�?-y����>�����ŀ�+��}1����8<(��Ajj��i$��u��^5��f�[*ߥFoh��ⰺ髦B�#ώ(j�Rʆ�M���gb�LZŝRQ��؋��$�[J��^�������g��B9S���]�����Ѱ�eMV�*Ƙ�a{E�Z��(|8sG�U� 6�BRď���w��l�OB���)e�?�5@�r��ӭ�SJ�c̙�s�0�����GUU���\�3kA`�\yi�������jH�A��4�ɍ�$��@V�_PF����b}��A�z��i��f�-�"�"+�3��
����!�>D-�4V��KGH��w'�W(C���)؍���u�+�:Oq0��}��c(�RhV��+����6t�iE@�{���a�:1�"h ��2_��1Q�-]=YN�*��"o;xd��q�m�(!O��S<��S:���ݭ�P�W���k��O��� �1��j�����-��n6���o�Q���_P\(z��}�@�4�.�H�''~ț��?�7�H�ΰpl���2�l �;�Ò<�w���T�A;2�+���Gh�E�(�T��X̂2���6�j��&���?�