XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\rQP�!�����Br�:L���R_pݠ�JY� 1i�/F�b%�X3M_��lX�`e�d&����.N���c���V��,^;"�Ҋ��b���J0�ē���V�z���I6J��2����,�A�G��^�_Pp���n�d�mOk���Z�-��W�Ѯ��2�����o��''���,'��xE���95��x���3a=|K�kX
۸�R������Q��I��.�It�kջ��I� X�|~��Ќ�3�%wQ��sc���z�BT��t(��-8�݉�.��6z�Y���~C��ID3�'��eX�?��Զ�ixv۫8>!'?M;���>���Yq�$��-���׎��u��qz(>�v�;�/9`S�q$�a&�x��� �Rw�S&ɵhkC/`�F(O4=��w���?��DWpm�Key('�!B�yG��(�B�j;Ry�GV�M�
�z�0����թ�y�Vߍ 1�9�l��ٵ���c��������zJ���Xw#m��$��|��fX��:��'��,�*������x�Z�7�aO&@aÙG"W�~�����C�;��(���4.��Vs�Ll���/P���k&�q��#�����Gd	q)�t}D9��!�[��JG��lJ�b
P�;��<i|��Y�/a��l��&�
%�y�×�ʹV`��F�� �plJo�	;�`����6^A���q;	Q<��h�{���
���=#֦j�$���XlxVHYEB    1cf5     790�,��9M!D����-�O�&+	�z�`�t���4�F�N j�{��)��7f��=H���Ve�IL{v���߭`��R��`�O��
�C�:���4\C�C�.O�^��4y.(hB�ި�j��*��DU�i�{(I#����r5�`A�=����M�V`����$5BmH2�G}�� �J��_D�j2��z@�e�ҫq�'��C��z{�����/��&��(2hP2`�PE�
�Z'>e��E�?}U��Y�G��/FH�E�43 _�<��ȃ ���/���.�Z�U+�6��V�rDo���"b�5�+��})�.J����/�d8=�K�Ȧ���㤂jx���9B0J�-����2Q8!�w�X>���Q9����,'�i��/l|	n�2��M�ekVa�,M~��s�N�Wl�6H��l#>����	�'�Q�*��z1�y��Uu�9����_�^B�{У�[Ge��h�n�1*��P���AG�\�*=���f0W�4k�$q�6ɣ�`���qB��B�֤%����b���n��⒫XM�C��B{� ~r,^��h�S-����h�3���ň�\��oǪ�N����n�o D uۻ�P����H	�0Q��y[�ډ�b=���!�y6���Y����C�;���Fg�@�U��U���x0E'M,���ƶ�p5�H�?���i�|]��%e���̠[>ǯ9�� ;2�L�^�v�to{���
'��j�� �)&2ѿ��NP�8t!�r�����biA���ۖy����{�t���ɲ�M�4����c�;��?f>C�_�ʖ1�$q&`��{[e��͕IL�=v�x���������V�X�ߕ ������#��`�������R^�7���Wԝ�y��J�jlU��H��z�6Q�!��5� �^#�E��Ǧ#�=/"�1ߴ���_y㲄<���?��x���[�� F#H�YhT�T�=����]ꩥ��*-���>ej ��9h�JǙ/�tGd��ʄ�p|Z�D���s�8u��P��������p����� 7Ws�9���D0X�$� UH�NKW�:j�?S��a�Nd��Յ7~4f~�d�����3�B��,�h<ƺB�C5uA�N�^h���v�VZQfp3�r��V�b����"�24�-}4�Q q�'/;���״���瓀5/�Y�l_S��i\�oG�2����@72���dӻ�ޯ<]�Z��b1��2�yXts�	�e *V��V�?d�ڞ|��=�����u�U#>ӫ�[��S��H�ꡭ
!����R �o
����%]�&��O��>�Q���F$�4>f;)D�;Z�)�8ݞ N6i�	ۍi���;�_q� Ȋ/.j7WD��r4��(��!ɪ�LV��3�9p��&��wrP���r��[�H �@��{�r	��]�%�T�]����h5���Zu��n^h}�ǲI�u���6���F�+�(.vM���5:�uZ��F��i��Fu���S�gF�h��#lyY~��$���0�S,� �?h��m|����ya�y�~�P��b	x�����[��^�s�o�S��x�@�.+�}}{��X@�	���M;\�����t�|�#��sK��'��ԋ;n	��.�!���,�o�]���x���me����;��7f�q��Z��4�D���W
i���{� ��64lؕ�������7�TH�ǀ��P㿜ӕ?��@_��Ƴ��$��I�_��4u&]5�����k���<j{�(�Z����mYv��Q�Ձ�Ss�ق
t=_Q��@�K�Ai�g�����)�8l{�/�(kՄ���v�����zR��բ-3�Sd����� �)Fd��h�=��Oi"`�˻�U�ǥ+H���Q�t�%��P�