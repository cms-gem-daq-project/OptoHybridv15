XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����xɁ�r[|ã@
٨�,�͑s�ū
��-�y�6�6��oCB�)��E�[Gڍ)8Hz��v6߭�Nf����_:��p,�~h?�#�0M�Uu��r��E�����JGy���Vԥ�ABD��k�2�B����ϭD�z��'�B�A=8ܙ;��9�=��iW��?��-Ǡ�w-�Dw̹���mX��7Lt�X���I!P��e�������������
8c�ܼ��#��4�����}W����]@����
R���$�)efC��`�I��J�O�e��0����|RJ`�S���Cx<S�B� 85����y���+����A�C�WC@��y���;tLY�N��D�4�)9$�b u���؎ko����ʋ��xN��x6�U牯�v�������<۶O��=�&��� @&*�=�̮���,�o p#�[�٥�,��N�|j�Hh[-� h9� �6OC4�FG'���ZA�5�����*���d���l�H��x����2�A���P���G;���E(�1�xGVp���g*�$������lk>�V�sa�{�{���U���mm��]ɰ�xJ�<eҥ��e�C �y7��H� ��k�u��4�J�I-K��_�zv(���ag�$+��k,��aĭ� �u��(�K��O�,ٖ2�������N������&�����4)�����f<o���J�l��b�*��dD�)�pg�M����J\�i�Hd6XlxVHYEB    1b22     760���rb�����Bv�ӥt��� 0�o�����2te����Q��!�3��K���^�x"*{7�a�R�͘��qX+���{�sbt�� �E���g��~\�\YP΍kC���֖B)�9,�x��zYc��;L����[
�G�$T����I7�������*!�U�pa	z�2�6������9�:0�Ɂ6m~�����IS�o1@?�ۘO���.��8�\o��񃌄����9IW;n��$���t�9�p�
�W�M����MH�5��qU�=���Ռ�I:�a��}�ˑ�C4~���^Q���Z$�d����D����!�Y�*�TBg{;��9j�9��B�W�a�=��<���g'��Fl*�,G�h���"�x�>4�C9i<ߴ��M[Wk`E��$<��w�3j��3�>��\�+���Dm���#���^q� b�7@p�I�j|�{��uҵ�������{�=�����CA��Y�nѦj��3~h �TC�!]��މs�qSo���v�fޟ춞�-�/��D��1s����̄[\%w�3�/�I �~������!�{L3n1���9%䏄Y=n��,?P\���&K836y �,4�����HP���)��(��z�Cn�ǚKaSrJ�\.�INtW��	��������2�j��S�C�I>�_������-��sAw���=�X/u7��D� ��,Z"���������B��E������8XgjN�2�t�P���f�Q���*�����ssG!JMɑ�N�8Z��"}��T�ƃ6%�Ҳ��<���H����s��A������'8����N�����"!t�X����$Kz�X��?���6-��o��U[h��Dh:Y*���uGuV���{���b2��`@*�����{��?k�(���N@K�&*�t��[������<Ά���B�=P+=>n���$�<��g�������Di��}��j� ,� ��(D�s�n<��+�")�u�E@ك���.�_$����/�h����8�t���˯M��
��k����:�a��	N���q��e�?��H�ec��;H�%�`�&��
����֠����
���-9+b��-yZ�������)2����1��
����6��-�_>�厑i��YS���C�c���TS,^��M�q^����}(��v9UX��ì��Yg��,Τ�������ԏ%��&1��ث��{���_���.\U���4�Y�CŎ�pZh�l��4��v̐�)*�ѥ�}vGL�_V͙,�P*���Jupz���:'�z?�T���<|��yw�����ݵ����"�$dޡk�bY(Blڠ�4D�.]=�X҆Q�i;O�ˀ�\A߿��-�m[��La���V�N?�� �g��䫧gᓺ�Hdގl�Ym;�!�	���m�3s��
6�oݯ����Ʃ���?��v	s��<h�Pź&�+��.N�|bN!޺X=kb��Q0�r	E�
 �Rl~e���߇��?h?e�vж^b�pl��ۀ�F\����Eن˨?.˨n��+n�/i6��; ��.�/eG����w�1n{��(�R#�7��6$h9���w��eN5��2l�N2̂bC�8bv�I��ћ�lݍb�sDר�����
��={F*�S!��o��
��n�n
e�W���|�M�6��?Q�tJ��L�{��w�ZkU�'fg
��@��O2D��ArT~2�Ju�<�ݛ��������^{r�fb��y���<�nr�{� ���\�t�H��b�"�~�7]���,j@p��a_ O�x��>��J7��k�c<��2�]��o�Pi��ѹ�<u�&�<�}��-?;��gKƬ�z�