XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���tPܧ���R%U+�X�?�6�]�c9���Z�}�.��f��c܇�y������$A���ZW����U�]!\u�kfÊ��\�9Q�b@+EHH�������!�.q���Zs��Y�_����>!\�A�h�K��ON�_jp�1;�$����&�è��&�C�M���|h�,�o5��S02Jѩ��l膪�D��>F��7<x�CN�G���*J=����
Qa%��8~Qv�E<���IG��7,VǢ���eR�{^�h�  3Q[�r����,��>�;��q
��aA�ǅ(�;�����]\`���O���Í$� Ek|��V���o�3��Nc��pQcH+=�G��ؒ�GǊ�R!P~jHm��7��&J���e�Y��).��C���� �O����B�O�'	��	t�B�tjG[ $�E��06���Uퟪ�����lV��`�a;Bx���P?	��/H�n[#�l=|4A{7�<boL:�Ы+�亱`���I�,��I�>��9�x�N-��P��E8b�
�y��ҶxP"��7�kl[��=��_ӟP}��]��1nZi�j� ��1��Tv��"dt����żt�ADd9)�1�7%��U/�~O1�t����q+,�V��S���;T:�q%K��#�Y�2��W>�����_�Hj��!=wE���y,	�$�B���`���G:�P��S���F):���N���N��]��NMH�k��<p	�"J�[g�{��$�B�XlxVHYEB    3248     930�t��3M+�ܭlh��I�!6	d��A\����;��*r���̺�A�-"]/�,[���D�I�R��jrM�ՁG!�T�+����P�2�kQ�q��
�M@L5R��ee�9��<N�*�J(�W�sw)�L.z�(K�6=aBY �R�}�qs�l�z���Oֽ��n���@����
*��RT�|�,֩	���o�#��r����Uҷ�HŏƇ V�����Y��tMi��?M�A�y*�T�rS��	m�D�m�@���ʽd�ź��;��*fl�+�R�"�W����_�B��s/�t4o�o:����/�Ł�H�C|���y��&��6t��TA��n���<���xT<N���V� ��|O��Pь�q���3F��Z1�SQ!�cQJ�`]�W_�.pv�_m I�p~��Œ��I��'����0\+���%�{���V�!�G�v�⎥/0W�&��FW�j#�7M�e�K���YM�6*�E۰�	�?$k:�X���a��}�&���z[,,Q��YAY��5Q~��1��17�2��'�e�M}`T�E��(�� �����h� rG�ɜ�{�>]��w{x 3�;E�xi�C8�r+�+}�[%.��Q|��o��R��w9�G&Z���������Q����.��O:����GC��d4��>Bǒt�����QU����E��@36rDD�9ʈQe}jۼ�!�tL4�<V;v��T`�G��2��+�u�]��N|�y���_2���)`�cD�q�v�FI �F}�2j��b7�"[��iBp��^"]V~�8�`
C";����]떆�[;��O8"�: ���+�Z����6�{�@��+a�[Y�2��l�`���Z|(̏Je��M���9�x'X�xX��w}tBX�}R%�� �AF�n¼�P��;mF�����7]��T�;;��@Ck'���$0���ٶH��#�%����~���:_��fi ׫� ֻ���=]ޫ��0����1��S>$.�t�h�o�Ϯ�a�;�U�� ���yq�px^�u�!��A��W[щDڂ�GSБ��a&ʀp�R����
'�DJ5o�4?G��a���2��L*����i9�C��:6:d�����%&�ނh,JMEN��0fPg8��[�,��r3�z���@�T~)�CT��ە�#�}g�S������0�u�
hgv�x�I��m����N"/	em��s��.D~nD�iE	�^%E0�l-�C%A�)oPg p��$]~�������:�>˜��=�d� �3N���u�������*�}�Oq�$����$WĮk���`f?���t��`��6���$�ʶ� �cK����@��3>th�E�Cև��5�} ���9N"�5ʅ����'�����F� ,�dD��Y�N$�%��؞�7�r9�wrzz�r�� ��`	��% aWEN�P���/�'Pt_eo,7'�Y2�m5wcH��@� ���U�[EZ�;��o�W������qq��A��S�H2DI��+7�'m��<��LE��-���Fж�/4��<���a9.�������D���hS��Z7��]�gw������쨡|�'����D�#O��?c+�e��G�E����L	���/�,���y'K�3����ـ�Qf�S "�]�1�f��`���ټH�=,Ҩ�}���t��'�S�,�W���UY<f����0S��8��ԧhvB�%v���
�×�PD)�<�?!1 �|{�;m�h�pP[��3��X:(��u+�?8���'�PN[�i��˥��D)�5��	&\����1�q��?x8�(�^�a,�~�ﾒK�eWL�c6���4��݀\&�^R[�>m��%J��Y5u
�Z��V��v���o�h��It��$�ȋo�&�'H����?H�����ٕ������50�̘,�8�����U�����|��eB��},�WG�~x٤C�.�|�.��T?��?��x|��U �z�d��-�^Z!�*�b
+���)4Bn��ڳ��IK�<#yWO�Ŕώe�c����ь����+����'�� ��#�R��s���6T���;ԕ������300��\N��X+�4�����$�u}����C�����jU����qU���fi�������9����+}�D_ ��}l�:��D����.�� 6�:�AW�;f��'T��;j����-ޒ{��y-d��wǻ�rL����%����[F��Wvht���!�oDG���n
��s8����1�}�?^iz`cB_�[�%@�.��Kq�S�=�*��a�kp@�Ps���S�