XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{)V�-<��j��A"W>ؙ2\�AD4��iJ3l�fb�S,��@�.�)��{�V$�8#�W�Y O�n���M/q�� ��C8�Y8/��,oj��h�ț�\�����w�Z^S����1
h�gi�~\⃛�㵨]��7!������Ϲv^����њ�;:&[&j3{4���s����r/��y�͟l�~1�9���O}�B�h�"��Vfi��x \&]��ˊ0��K�!JƼU�C�UsGH`���aZ6`�J��C��ȼ�ڀ�~m�r�����~[�}���g���8i�JljC�����p�x�]�=�+9�e��L;Qf��t�5��Q��0��l�ХC:�;B�6�P�jPU�{�+z��`�`�J
$X��/vF]�a���A�ۉ�J<l�j����$�Xm���t=�*"�|�'�lu+o�˹��`I���kK�+J�́�U��ra�_@��!�!��;������t#u�,Ro���� m����f X��^O7�4R��3Ӏ���lihe$�(����v����Nes:#�O>衂��л��S��[������O%C/*�",�G� ?Ll��p�ul�`.Gc��N����_���͌3�=@���]�]L�[+p�P|r�-%���"���
�ˎ����a60��|���1�]S�Uǡ|�Y'/��;����? M���_"�'9��|�X6�k��{1�{"�?D��}HT�d�9/F��N��1*�Ч6ɰ%�VG��W�ʹGX�C��|�*y%T[S�XlxVHYEB    2863     8d0-{5�@R+���^EN>ך�ю\qg�ҥ/�Þ��~�<���?PET��4.�f����4��3l��=ܛWǔZf��wg�k�0���=;Q%���b���JR��f��?0�PBp�V��<���ApR�\��9�x�o`�ϼW̅6�~6%2{W�����t�)�T��e�zd�A������r�L!ĊES]\�uz|�Vyx��$ߝP�><�ok��֪+����b ���V�&�e��U��}����m�l�4��oQk����=���RUqp�:$�A��*yє1FV���#�5	J2ߜ0��]�"��D��I������ (t'�~�����������=����2�XDZ�<������{�e��;ރ�j��<	����/Cjq��E�qî���U���un4�6��nl��,9f�7C_�Io�yVm�����UN)��f��˼ܓ�9���S33�N���� ���ǧj��_�k���̴�@��0!Qm��W�z�O8;K�H���q��|��i��"�Ē�{&�:���p��e�Ji#��U9��J�����(&"yb%,�8��?�i��*�}���43F:P
#}~r�·(�RO#�נsX���V���.�"w���
�{�VYL�l��D��X8�le�{(�+9{��jUm6z�P~��Z����g*3$	������VWr���[7�f��P�o��5[��j�9��/��}@V�c�
�0�����-!���JC��џ��"��ּb&��vv���w�,�-���].{�|��b�,�&Di��ݾ���4��9��F�qSM}��	M�򊜎ʡ���W�:�?8�#�����bp�3��*A��,�E�섟f�Qytn]�����Dk4O�����dh�5�Jlzmm�?Ͱ���x7���?|)��0ڿ��TH�\6��F{�dU=�аBL*~)�n�e����8��࣫m?,I"��}s��6POX}<QMω�.���a-&�Fv]�i��q����tx�d����v��B�Z�v�҃.��û�V�8�5�VEb�e�����2k �uD놭s�WU�<Q�]��^p O��<�&��z Q��φ���4�v^_�>"p'���0mĂ�����~��!_��s�Oׅd���=J����В��u<����#y��B�u�[X�r�}������c�s:5_�_,��7xZ�(Ș=O�H� |Έ�y��(`�/�
���n`�d	�\�J�r,��ꌣ-�qt��1�4�ø�l��q���!Bـu#�����Qq��m������K9�T�z��~dT�>�Cs��Oݼ@C'�S�3vӰc�}G���
�Fks���;�I�6�N�Q��y!��E�v�P-��a�EH��L1�v:W`�(Ɏ
n�H5<SD�������]2gֱ�؟/ G�o����0�,�/CS��zjro�~ԫF�_����KX��Br��w[b?�7�O� Z݁W����?"��V�~Dʩ�['C�q�$���4����b�$�,f�U�毅��B���k{��s,��l��N��}����BC䌣m@�S��#hr�?��Z��*���-~i�UmgU���E!&��iA�%@g9c�C9��4h�X̥S����p֯@����O��4h�s�oBy���q>5��he��t�>E��i�.b�x�(����BJPk����.,����L���6�SznA)=��	�/��p!py�q_�H֑��YI�n���L���H�Z�u�|(GU�#/Ո��	ibhY?������}aaj�AĻ��L��`^�%��o�!�dT�S?]k��$����l1G�R/a/@X�V	�C�l� �ءt�ٻk���)/.4́�tdhA}ҜQ'_�������0�3�������ѡ'7�3j?�t��6�����̭V7�ҝÏ�Co�tx8�,F�6;S���'�����)tP����O.��a�%����m������$h��/��7��X�\)����8:�yB�6��'�p	���P2wO�;���87E�~ȗT��|}5������ᶈj*����h rR5�BU�>��i�0c�|�KHLl�^3��C6�+D=�>�Gn���G����-��Ss�}�8���LLʵ8]3£K�O�bT�|T��f��3�US ��A�;���� ԁ�A�J��N�n ��va�k�p��B�� Y