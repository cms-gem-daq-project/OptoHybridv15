XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?ʱ4zk��. ݐ'�>%w^lI�9�ߊ'3�%Ԙ/�@�2�K�*t�'\b0&�8��\��.njc�vO�� ���7f����5�<��U���T�x���=�ۂAf�z���]�wF]��rN$�6�篛�E6FVͯ�2�?��a�4�}��S���I�0�M�����%�t�є3� �)�V4�����sp8e��l�m�D��M��í����~�&�BB�QI�̭�lu���#6�SwZ��dj�?b� �L���B��۟�\υ�q�k)�����������@M����V�(y�����C�� �á��1g�k<6eü��i��/���g>$y�8[�T��l|^���|G�΀��z�`���Z��i�FךT�i�>�b�ѿ��`�U�GP�Ỵ�~%vY��C"�3���]���^�� S	Gw6�I")���ѝ���'JP�n��޵�RO�\ґR�����&��$�ձ�Ga݊�Q+4�d�����}�>�%~]qW�%�,3�yE�����b�a�/���ف�:oE��b�%���E�R�b�:b=��F��X����������]7
?��Ƙ��g��+Ǩ"���n�N	���;���A*7s)Fu���sO�e�u�7�M}b��P��}�ϗK�������V�$g��/���(j��t�r��l
�������L�����j��m�4�>�Q����ѣ�(�+��-yv5��v/*�#m ��4v����M��\�b� F�,y�
�~	P�:/���LXlxVHYEB    88a6     d60�L[����Cb&�s zA{��0L�T�H�"w��~�;�H��)R����y�f�
],ht���N�����mÕ�I%��U��A�Κб��lX	­p�5Ϫ�_U�K%j6��ić	Gߺ1��B���_���+c>��~��Ș*��(Tj����"�s�(p�#��˧�>�y�`0��j��ՑP��p{�0Vyt���3��R�������p�R�s)^C	]]/���;@b7�o�s�	Ė4���⒜Ec8����Q�ő)n����1��W����/
���>��u��9x0�,�w"a���t���:[����𜒖a��M�����q���?��A����k9�y~Q��nSWq+,���Q9=?�O��w�{�u4�^��7⩁�>r�VA}�L&�����[^c�|�oW��U��:�Ο�X$��0�Ыw�^c�� �®v�?� �]�}Z�� 4@�?�!��T��΍�E���庖ʀ�q|��k�8p�&L�pȴ��P�45~�]�X{m#:g�đ쒥�i�q�<�e ;N��=3?E��=����I~�M���#8_'�m�G�eV���
HPg;g@�d����#>�^h��¼S��ޟ���$T~����X?'s�+?�6Ažܡ��~�hOxVM!=`�����$x�<��n<u��p����t֮��H��C���l�/��T�*sYpx��ݛ�J�oJ�c�q8��G�N�R�((��-
z׌^��oʅe��Ĵ�����i�������ޠ��e������L.l�nJ[k��^b���7�pS&��J�E-v`�Vu;��Z�m2�3�ԯa�OL����'Q�����^��z�ߚ�s{r�����x4����K1$z�?��jn�-�����φ�NY���g�V�\���%#��ڬ��!��V@M���a�h�R��l^�)UZ���`�s����Z��E*�	�vy�2�Ҵ�1���5����V��h ,pnҳ��1g�A'-��zq?�J)��=�C���i�*sB�Ij�.��m��ldalU�b��^Y2Na7�[����{���q��"��� ��krL�2_'(�-N�v3�~�a2|6�Bٓi-V�RwRٹ��f���6�D<Y�.1�s��Y��ؼ:mQ�K��OQ�B�yy�BQ�]>�
�#Rt��u$\�Oj��V�����W�_UT;B�+C3W�-9D�Rl���P�����>S_��|f���ƶ��#347��n�TRjF��o^�jG��6�L�D86�C����8&uǷ��nΜܗ���3.=8��?��4�Q.Ԟ*~�{_�u�yIo��η���?�=��H2tɤ�kD����'H��"&������;�T;Z����'�x����"�X@1�9��;rЦ⬏Y��e9Jd���N՗�{��ҭb�^�o��w�A�y<w	 �o*��l�5� ��	4j�ZN[�嘖��Դ^U�C�Y���h�#��z��v;/`��t�D<&¢����/夵�\����.�ha~n�Y0�eY��}�&�p�n�=Φd�0DUjV�^CT�c_w~$�O<� �[��&��^F�\��#9f
��hBԿ$l�"bݹu��&�TIM(x*�n;�t�'��xZTu��@�X�;�GP�@���uK��}���>��Z���*LMOZ911XvT��k�HƄj3~���9�6x�K��h�;�@�y��V�e�#��M�+��cKp/���^R��U����4z	٨ʹL��q���w�kD6��~b�o7B����5z��#�ռU�URq{o	�ap���|���I��<u�hMgSXz-�g4Qz���a����_�f��l�ȅ�U��\��fѰ��ϣ���������$�2��컁r���8D�CI��}�}^bv}پ���	4��1�Nֳ{���~п	\�1�����W�q�TRR��!�>6�b��+�?j�'�r��i�	;�c7�޸�����%X�������-���\��t��'����	|"�4�x�u�����H�(Rj���� w�ܔ�¦��@��G6d"o(�c������6��S���J0Z��������m�o_ӑK�K���ikݯ�tů�[�s5��?�����dH��b�:D[{���F�!Iw�V��Y�+����O���_���S1�n�GQgX]��~����@�OzF�p9X�'۳�g%c�����.��Gߎ���vs�%�y0��V:F�����+Ѧ�2V�h���V��~H�T�S-�M�pwDHA��	!A}_��|U�1�t�$�yhV���d�!I7�|d+�`��%�?r��  d�f�����r�7���
�hϹ7V�-�ͤ�8��$�[�����P��\��vv,x�k�:����+�\^���;�qC�o|��B���w�#jإ�v�:'�#�bz�J𐺍�V�i������%�db�L����f���z�P���8�*�F�zǘWU�t����V��"�'n��S��?�
W?�R����LFO�^�A�^6��dcT1�I�Ɗc#%��ʀ��v��nk~�l͢K��lHVХ�pNX�k�n*�h�v�J:�f+.۱��3���d�����OJ"�&��2�[t�~iӫ���P(����\�x(Xc�D���Û:>��|m�A+ ���ۗZ�=��A�w��O)��&\TN��,��0����g�9�i�H��ê��MIgU�b��S?0� ��l�Ø�!���t�� 3��D�UF�7��g�w�!�.�x�5У��iv흺@nf����B��	`�q��������{'N�9~[J��bA]H3��tP��s�0���A�r�, S�����9�5��^��8MV�Ca��	�l��y�Z�	���ɦ�d�`�eR�;S�b�v��,��ı=�%�q��\g�vt�
�"�7����*=ܧ6�� ,���~�ӝ�m��h�9w��r����X�d�P�w�X�@V`�r1�~�ߛ�nx�� �Ø��o/~2�M��m��`a��D%��I��g3把��~�qłƻ��2b�]�l�����11��w�B7ǃo�B�`�!UGM͗���:�2[���<:O(ƾ�,q�a�q�����Y��xY>��e{q�s\7�v�]@��~�{�,��uE�q>�>�d�F	$'$��,�Hc��*��5�>g�,��}�i�$��[�9�4�{��y�ÿ��
�TH��m��lr���Ѡ��G��7����=T#�%%��=	'��_\�U��ʍ�*>��@���?��q
��o\TJ�銞&����5�5�2L��:?d�K�p�K���*@�6�S�	��� ;��]j�80�