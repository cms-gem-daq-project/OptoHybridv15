XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����<��^v�L>�����𻎡3�aO��V�Uܢ�J�$o�O�R$���� �a&Q��Kc��8�l_��B��<�����8�A
����BW��-ׯ�`P���Ys�!��it��u�qJ.lLa �����|�`��-�]x>�j�>g����V`N	�����n��Շs`��4Yl�-?�x���Q����-�>�9�� U��AI�$��v��#�Q]!f*�R��@Հ{*"���HB����+ݤ�}_3�8=� '�!�&�˶9Z0���~�)nV�pi�,����������T���#0��m�����73w��Gl�,�}"eUޫ1�F�')`��T�xAg������G b)[�˚ߺ�Z�PF܏��Sf�bbM.�^z��M�$�a��	�%m��omhTD�Ւ�?sn(���\��X�)�	�H�K0�����Yt���֫r�|��3l:2���½S@��mz��I�U�� �mX��rNhߟ�F�o�,T���H{����a������Ʒu��n}�� ��"/���F����"�L�'�^P[��g�2����[��N/�����)��{�n⇼^'�����v�T��(	j�����e(� �l�ݑh��8�����F`X�
��؋E�DE;�,3�d��<�\+r���7a�_�+��"V��L��L-�)l:Ar�)��!Nغ�_�1�QO����O,H}�;R�v�� �+5��^1/D�h.�8R�Z�U�Aj����Y�L`�����흩����!XlxVHYEB     a7c     440�v�����#��ܢ��%B��`ޑ�Xu�̼	���]90ih#;�"Y�O�ł����F�t�y�<Z���L8��webr;�(�>C�
}9	B���U�n������0:x�0!�Qܩ����L��G�QW����ʒ��1��	��R8�֫X�X����#�z��&�1R",9���{��쐟F��i.���o���/�m������.���`��[#��b���-G��S1����Y\x n�l��?'cg�U�?�ۇlj![غ�!�gڟ]%	�1��2�Ш�eC��%.s���f�P����!��N��C�t�)��70B|�F'Y:��A�`��Յ�t-�nUGu]RQ110�op��hr]1�������g�/�y��I2�cX��uX�rr��<ٞP�z��N1
�ka�G������c���]E����4�ȓ~#rT�|��99��5�tI����l��$�FS^�h���[ח"y�A8�h�5�c:�y�A��bU�Ė�,�|���\�K�AҖ{VT����xh���6U��v����hv ��z_7m�2��)�j�+���5�	�Ǳ	��5B&qKڙdy����U�0�`�k� XD��3҈x�TԊЌ�`g(�����"8��	+���a�m�W��!���\�%�#�	2j��KU���?��dK� ��E��e/��3�si����V��dϩ�:��p�/��gxu&N)�<L��L��DW=%7�+�8e��mH Z�y����~��PN����"B��i�A�h�h�\�g=~�) ���8�>|�}�@�V��w�a͆�%1���l��GaH�s]% ��;�E�MxM~�{��[�p�녋�F)]�0+J��'E�{n���Z�5z���|ʀ��4_Ⱦ԰�$;|��v�M�4��'�ͷ����u��E�
a����x��$��Ь�O��5 )�Vck�f���fhB>3k4��Ck�D��/X��,�N'����r;��Կi������֚���������k�ہ�+F��(M����A�S���P�ظ�˾�a�:�l�Pua�o��l�r�|�-��Ǻ��#�� (