XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g����\���;���ZY���E���F�X�O�T`)e���n:��8q����Rg\���a�ˎF��/y3O��"yZ��GQa�#}Sf� 8�
�� ���g���<CV��.Nfq�
:�H��|���0T�� @�`s�L��X�90NK���q�~��d���b-6\�@�)��D]98 3N�2�R�c�2<��.�!8}K^'މY�����S �vl��c�G��^�����[v<F���tϲh��,�n�#q'i����f!C�ng���2�4X�iu�%<�>u.ӑZr���<��Rr�:�*��LE %v�5�F�dtjY+e�{���Y=���rHw=^��ś]ϛ���&��>�W��'V��z����h(����bK���r�|L%4 ��ZA��e�H]��
}{��ݍ���Fy���U�j(�ʻ{�2��6�P���@_����[谂_���aU�S0׃��8���h��r���[��R���),�;<�s8�$�>�??�Z�ق��q�=)��K�ft5:�Z0��,��(�N_�CkA��U���5��z� �f�^��l��i,'1�e�����=9O�4�tl���=]_��Pm���O^��2�^6тg�@ �np�f'��x�o$>�/K�p����|U>'���K��渠L8��Ir1s*�k9E�g��c��U�~*���%�*���cTgE;�=��i"��r��8�{��t�p�_׸�;B������{D��rF�XlxVHYEB    1621     410W�+�zM�!_"�+� �B *����P�XR��+�Aᰈ�q�lQ+�[;�oNZ��+adyƛ#Y>��&�)u.�p_W���$���Dg�Ux)�bK��	O@P�B��p�x'@��ho�{�Q�a��r
� �CI6c'Z��6�\����>�j��� �c�p�����g��V�{:O���r�c!S�N+�u �-��s��7*Q�� ��?Ѥ8fwpP����׹�'B�&������G�_�-��6�*ַ�:��#+����K�T=~�M���q�pp &X���Q�D�<��M1��4�р��x�}�<�3<�qgk�=�`�b���T	u��_��UsS�z�0�;	���|:���]3�8f��9�M�{F.��v�M��6����Z��ő7�����#m.��b�)v�gNrP`xl�j�\a�l��̇o`����[��!��2'�����7���~���P�$��45վp�C0*+d^����KYt��Ś�~[b��K�Ed��#��.T5>��z�L�!Wꐠv�8�5~۲̰>�����=}���A`�����%���"AO�O����,]�J�ܻic��DJ{'�	�3�x�]Мˏ���E~M���}ȗ�89}xw�4��y����;K[�as�/O]�Ժ{��'������l�j�,Q	00ۨ��&cT�0_��	QI������;����}Z�D,۔��i�U��~S��.���������J
�I=^:Yx��n�?w˿�ws�-!�1��*��@ 2�@~ij��k�$A��P�Y��$i$7�W�y6+�e�(��F��K�C��=M�ʮ\��G�b��}ԌT�;n>k'�)�.�<uE�~�
���I�(B��,}wTf�'�P�Yk��Ȁ�kKz����������ST"��rAh������Vw����um������P�)V�~�8�L�3�M�ݶ"��2���Tl�o�@�	�џ�pvt�(S� ��񗴢x�k�ge]	x��B�!�nr�