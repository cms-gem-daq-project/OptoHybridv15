XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������;���} ⭾��9�0����1��G�q��9�2���ٗjJRQ)ch,8Z�ٍ��f�[(Hi	 �d����Ԃ\م���\vׄ�|y�h�)�ܵg�,��(����Գ�9���|INf[4̥��(o:�M8����ѩ����g��?�c��O�,ك�07&Y+�K���VP��B\L���l� ?�ޠa�C̽�i��t��O,����0���Μr�3~
�;�S��)Z�ݹNt��aTm��q^��o��#P�$%����� *?�_4��J���b>�`+;��Q^/��Rn��+;��${���7t�� ���mU�bdq]l������Pn���1ޢ��HՌ�+�a(7\;�*�����g�'��wV�{����ݤIh2jv�="�:���d\��Ť���iȩ���`�e�@X���R {�0��J1���k5������5`�>��2^��"8�H��c�X L�b��̍�|߃�6P=p7-|-�w�r���cO�������^��I/֩����T?C_F�Q�g���B����Z]��y ?�6k�쪈��"7�x��%;��bx�����j TB04�bv��i|��=a����z,��BS�M1��P���������|���j� �R7	/E���r�p�|�Y4����r�����4�e z��ҖCKg�+z9�L
���p'���5 <�!���8vt�)@��P�l����EQS�˽����ű��h���Dy�C�JJ��XlxVHYEB    216e     8e0��jcA2���|PL�h���b�,�G���%�s��n�pb�Ņ��@���;`��o��t���_��9|/`�b;�Ҵe��Sdu]2:$G�;�ܝ����`����j��2ل��J��Z`RY2�a	>����QA���d��Τv�w6�յW-���⯧~}�HHYI�Ί�q}�j����%�9n�E�`KX�	�5`�=��­$���˛Y<'������f>=���>y����3�W���Kl�I�QmH��y��t�(�ڭǎI*-��U��'En|^��*���7q��dh�f9�;P����~3X~�6���}�\�Z.�	���3�?+�0��v@Xy6�%Y�|��[7���{բC� �n��Į��fDKT��z��O��e��=���G��rc�N���d9z"@z�(4!DE{����K����!?�3G���m�#'�=E`?��T~7���Θ�[��$��#@~�͋|��sEА3�@�q���0T��LqX_����t�P�4�r�b�j��qxX�	y����������*��e��}�@�;�*[`�U)�U�y�Q;���?���&��=�k��-4�+�e�|�N��3+�֪�>N����!s3q8�^���N9=sY��FG�����t����rFdA���Q ��*�i�Ԭ�A`�h;_S��bT7���V
�=䩞�6�e�ye�/>�Ba�_23���U��k^���$F�ܼe1nx�S�(���v�I~�)�X���Xٮ�~YJ��˹4���7V~�m���h��8iq���}>9S��U[/�	"Ǘ��J�m^��2�!�*Ck J����	�_0r��1g����U�|��8��mD�T�e~d	�Wf;��ԋ��`�>[ ̅ �$�.��2f��Є����U6D�Ԉ�c�AI�s��d�Qgw'tW���{gL�$�Y���4�z��`4g�æ� ��Z�>�mq�p!������R��`�"�~t2�#��b����l��}y��l�h��U���t���Y�sإ��T)�U���t��Ԥ���*tu�Ge�����f�\��2��)ξ)ȝ�e�P>�9��
�����b��2�]�
���s�C�7%�(��k95PV��T�D�/k��č��[}��,��k�҃�w�V��t�~�Q�/[��5�]�!t@ƞp�É_yky�Lӌ��}� ~�l���h)���S7&����Yu�����y�%ku��!�
���69�e*F52�~�s׻��dF}�@������K=R\Dr�qL�S��v�=�}��1��ւ�$J��t���������,��40~ <����!pq ����	��� 7qL9�(�H	���N��v�瓲�i�Z�Z��<�/��!�1�)�0/^�.VB�z<��ŷ���+��ۣI�r7¡(����-�VfX�Ŧe ��A����ډ���q��e7�bV�mn�/��)�w_k�d���46��wfѳ��^��Y�X�a!��7Y���F�Fq��X)�,�p�I��k���:AG%����}X�¢�n��c�gvu��t P�qF��=�g�.�
A�&TE(";�Aӡ�e�x�A�r���s�<���M�5A����~��l�[t����_"dv��)ի�7�oZ^ZH�h:y/_�it�-Z4�UgD��{_�ؔ����@� � U�+�9�J�&��脏�TcЖ�I�'%�C�L&�ZG҆-�p�X�k@��-����L������5Z��J�2�u`�@SJX$�|�g�rj�x?!y,	��$w�Aͤ�5Q�`�/w��mhj�����r0��&T�Iv>!���a,Xn�+P}%$���;�	�+qt���*������T�ȿ����ft�~l��0�]A��={ITyh��2J�O��N#Oٙڻ8�7ko�B��f)������W�+_����l�99X��S�������#�M�mHvEI�X�5�y��/怼M���i:۳�s�7 _G:�o�`�0,[�dif
4�1;��x��V�җ�+n$`P'|�t��h�'��O#Uc��m"�J��m]	�mu�.}�k䙨I�&�������WHM��1*"�9�Ӽ
���s�� T4���ɚ�j�œ���^�fX�3GhĪ���1^��������XLP�j�Nd�}Z$�}ty"��H�y�����%���}4�J�!lǩ!�O���l� ��
�'܉���
�u���-��(N��� {�K���1��G