XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�/����&�?����<��6/
��Ck7���J�Θb}��+���b��j �
��U)��1|k�ۣ���(3����G��y��T-�&�H.<Խ�����k�a�w��Τ��SA��'eƪdұ9�2��F��ǜt_pW�t]~�
���.���r���ܶld�>���Q� �n�*�l��&H��,����4�c �u�_@u-ʅɵ�"�}��_&��4��>B�Olc#�%'p�%�q��\$�j��C$+�1��_��Kg`?G����O7���y�R+yRS'0PXo��A��0o�&-L�t@���o|_
M)ſ=b�l$k�mR��o�>�U��̵���xh:�'gu7`�AIv�
�����=V��Cr���7��{��7C��!Q4�T��+ۻYJrT	X�>�E*=��F�h�Y�5�)s[��d��� � Q��O����i�}r[��SeI���p�]�en�9�l�pP��%^d2�C�R���ܩ�Z����g�Ǵ?��18�ʋ4��!t��X���!��(�U(��Ȋ������JT�En�ԋ�thS��G�<q'kĒ
���]�d����i�w���ax���l	��2)�`ZkA�B�Q%����1'X�Z�T[��Ř�k���=����7o꾷��%�'`����A�j� v�������Ze�-�'�q�֣�p5HX�3eݽ�3�a, "�=�����ޭ���4�Rrz�ho˓~�)^��`۴�Rᇬ��ڋ'^����/�aXlxVHYEB    7945     7a0�r���[jc���� 8z���G���{�a4�g첌V)�OU��*���<9d�!�|ZG�uV�ȴ����=�������'��~0Ü�jЭR=�uK]5�g��:`��QDe�qL`�!��D���]�~��Wp�\�|�eu�R(�z>�wH�����%5Z⼗�1��'N4h��T�����DK�}����g�~Lg�w�W�[�� 
§lN$��kg��n��𖂤�B�R����@ :k}���))~��4��H��U���\y�G�r�"FV�a'4�*�Т'~����b�9���?��I�1����F���}�\[�F��L�ʕ�v��ˤ2*O����J��2��s$Gc;w(o���\mUyY����Dw��l�Lj��S4Q.g�d���|�\���i\�!�%���vsye��j��.�z�Q���tmH{YE9�<g�͏?�&4<�\�O��Ȯ9~з�>T�������B�^d�#�3�yb�`�^!Q�d�����^G,��2*5pE?�W8�{��L�g�N�V`E����u�R�vyP�߲P�uҝrԗ-iE4��UE/�w�]jv��.������8h��F��
){����|��ܭ~~4ZF��-�9�N _pϯ��^�d���� �6]����؜�D"T��ѣ�E�z���?M��O��eX^�p��t.s 1��6��<��cq%�<��)�m(��Q��L�(�0j�����:�g�0!(��=��M}w�Mc=*�q��f�"��}T�ߴ���t	���������,Wt
5������xI�(���뙪���΋yo۲�f,��+��MY�C�%̝���NK���?1�{d:��r��� �@lIUC�<qTv)���L�C�p�aT2���$q��S�3z@������ͺ]Q�T�x9e�v	�n����G9��yQ����	���}
(4u�f��&�ʌ�O���A,��a�H#���Üޅ��>AE���l$�f��!M��iL�2N�
i�X_�}�qf(_gd�m��|���uЏ!���1N�w�<,ܵ3�k�XN�3�H�="D2LްaU����p�� �/ ���[�/�Z.6+@�.+'�e�T=���W́��b�T�iN����A�j8�Y{{7f2���K�X	7�}5/B�r,��rU�����S��+z2��Tx���v��Ө�?Տ�D���HD�?tT��:�Ϛ�h���v1/W<v���!t��U=�~���@(�=����x���4� y�J�r�ԃ��F���G����ؐ鲆�t�J�0Ǒ��}���P�z{A�'3 �3��m��s\����+�0��7����o�^*m�Աi���:"p#<��Q�Ij>o��q6T,��`���}�ƥ�������5f��7�O>����9"�����E\:-�vgs6�2�2����#es_����������N_�l�9̨(Ze������$7'-
�>�-9��jl�\�Y��L�����,���~�{j��9oqZ#դ�̪7�n�E��6��T������p�z���׬X��_�;�),Zv����=5>�o���"gvr���v6MT-�zh�v�\������ʘ&�>I��Yd��D��1�eF���Y]�g���
0�H`����k��]�e9Qc~���0�J���wP�7(�V�ɴ�s�	T�t��v���,����]�Ʋ:�4��&\�Q ɮJ�ɼ��ĳ�/}�H����;�%���.�.F<T)����x��&�$^�S�Za�J�}�qJ�B�B��Ԋ軁m��]�-��Ȃ6�m�%���Ӊ���az~cu#o=���5�"SL��.�i�8E�^7������*(������b|$h�0!�_�m��1��������w�y�2K�6Ғ�=O2ݽrp��o��