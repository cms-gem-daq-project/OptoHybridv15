XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6_+�
T�ġ2�6G�D��vM�Պ��~KOT��L���@W ��f��e�I�Ū��B9pCy���-�;�6�'�軭t.�8}C���Ld��p�4��;ˇ�����U�֞�l�yc�gG��/������BQ � ����)�~D�\�#���wp_�����x�U9���k:X3gyO�H���E�t:����)c'��F-hT*e�����r�!jIÿt�P.��E�i��_��	7\Gx�gT�Ȟ�-��L��0a��U�хmR�Jg�_�qܷ�g������&�jF�S�+��0����+�q
�U�`�4��!�y����eP�!.��ߵ�G���q��Tf
��A�:�-ХT��ar�uZ�)�� �s@���
�~��v3�3lO((3��1V�� ��ߞb�0�'���H!�?�-}=UjR:|c	����4'�-٠:T�������@��8'_�g-�#%�#u�FSM3�.�E��}��1h����a�ޅM
*Ƅ[�=c6 ����!7�}7�A��;_�:@�6��@����̈��,��Aw�|�^�q	����+l#�'?��"J~�i�%|��+�:�&��������R��eA?���mV�QO�ߥR���)�k�j��q��w/"Y}ֿ��)��(i�����ƣ�2�{t���	��e�u �)U�k���������S���� E�؀x���b�*&�'��eN]z����7��&�jM��+B�ߎ�'��E.������K-MzXlxVHYEB    1d4f     7b0S����#J����W{ȥ w�X��WV}���S�j���|�}��o_z�t���b9�&T��9P���]c��OJ�+_�M�/h�����zf���T�1ȱg.S���JX41���G!�*��8
Sp/כ��򭿍C��.U���	����ֿg3Z��qU5$�q���u-�u�Y�6�0K��:������v���_�|B���Ak
�.7�e��\��*����ծG�En������Y�̲\}�hH���:��0��8���&´|�����yQ���A3�j�b��1-�Y�9�#��T�-&@>N����~[c�1�d��c�?[6V�˾��h�;oN�nX(�����Eڶ\�,�ҫs:��A=�d��]Y�*/�Z�����bt��'��s�f�:ԅ�ef��5Q A�^��^U�̗o��m�Ł�e ����R���%}�0�CG�����L	�e�o�k	�/�=�6��V���O�|S�$7����.�3)��bKf�p�Т�\)z�IPl�?�B9�@ٯ�Ȥ:x���V�����΁j���=���}��)�Ez5�h��ۍ�a'��� �ͽ�>���I�
��&�#����{h��`�{�V�;���%�[��=��z�(d����$����X��G�~��'� �z@/Nr��d��bR֢�=�G�[-מ�`���g��ckCP �x�k����Í����
��gk/��V�\�V�Df����Q�r�/��r�wJ�ᴀ�kR���\�v-y��^��f�<;�S���Ǔ5�X����@���aʑm���Ɲ{�j/�8#����fo-^���H3�+�-~\�I��f}f#�0��򯙇�X�|��@%H̪����OFy���?���!%t[^��4j��
��5�:��x������u{>�Ba�Wؽ?�k���>��PZ1aI{��u�e����J��s��c��dX���(�*Ŕe�u�Ϋ����T٢.��d�/������C:{�2�o�\<�FH��L ��z�A)*�v�q�WX���+
����X]s�R^*H|�bKy��.���9%�d���reHV�@8�i�/�~ߛպ,%�KEÎ��P���VA�v�c�~kv��m^悥q,2��^"��}���z^�z�y55�sx�����3b����M5H��P~�z���ؙ8e�gj��T�z%�����R�R���~Ч�ӭ��@s�����������i257�^�ϲeJ��m�5��]W��u�Q6o��
\Û��l<0X��4�V�פM��.
�]��T�����c���B$�^x�OڤSH�DV@;U�}#��T/Q����:rvi+�r���B�yl{�T�Y}����4���0�l�u�~�(�zT�]�|1p|"]B1���;kd��D�Hm�l�;���)�D��)�،��3]Hd��b_Jx�.�]��j��ʐ �i�,�}d���&'8�BZ��@�%o�3�����]K4�9ƟQ��,:Q"l~�,f�L)j-�{y8Xn��=k2�4���q��Ž�h���2d�&��*1�����t�	VU�#��_��1�s�푍�ȥA�`a��T=���#7���Sq����O�f�ĸ��`�}ijMx,�c.b�f���{�<��U��\ӽW�; ۓ�.�S�7�v��N�>�.
��O!�L��,�o|c�{-�Ii���:?9��[���	��8�/�+]�!~��f���qV��ei�qs�jOտ
 �{�zR>���@�5;"��2��;�&�
�z�WuEYd�Q�I����e΃!l�&��m�&��t���i\�|�Z�R1l>?*�gWi=�G}�rc\�#)�4��c[@�>YJ�x�p�,�R֘qQ��*>����\y.,�.r�l.o�!��Q,[�Tr;�ӄNT�xa�[�����Xu�r�]T��k�ftҶ�d�h���:�`���"�