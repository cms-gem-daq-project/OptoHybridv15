XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����0Qu^�N0��|��ZAp*Hۏ]����tۺf�M���'N*�I�i�����y�$�bG��5|B:�'�	3����p�-%#^�V}°C����"R^j/��)uDj�F�	�$�?�����������)�)��_@
~�@'!����DF�˂^�B�25�����M�m���?�� ^90��I���j�i%me��[�[
_J'i(V�����QK�D�v�qM�?���i�#��j'SIut��)�d@���/��l6��F�.kbkbh�J�!��I�5|�$P�n������RZ�! Y��/���tx��T�X�+��(CN{�W=������0���ԅ#W�i+{(w���Rq@6:Ȁ�%��J�~3T��j�۶`NxukB�S.~9yT�7�����+b�Vlj�c�<͢X��	U�_�yAP*ȄY&���eUU����)d�خ���^���Kn���Y�n�Ȍ�he��Mّ����q{�DԐj������RMш�n��%U7t%�Θ{1��g�����SK����%o��=M�y��߇k��{߶<�6%e��U���N1�I�=iĦ�;��'�qf]*�����z�R�>7
��{8�L/M&�xסB���7޾�K��qp�+���kV��*��������y�"x��n�02h�:�Q�]�} �)2�0���Z7d6����ᇃ����0�tu|�v+���Y=�_�x��Gp�����_H���4$��W�]����XlxVHYEB    1cf8     790'e
qć,d�]�l��R�V�y�"̝���}�CrҹDa�z�ƪ�~W7�F��LZ�^!�(ݧJ0����X�S"���s&�B�S�ŕM�~3�N�)�� >(�3���g)17�8LE�1M�ǉx�TU6o��A�i[��ѧ����>�]�@S$��yi_�li�-�@�˫#�=7'%��0���Y1#��]��]������O��8��m����g,�% ��O�rC���
�.q��'')\�#|f��.T�eߵ��S��x_x�7��a��G�|�t�IqU�����2:�Y�f���)���
�F�@?=X#�*ҕ��V��k�J�yT�A���$ԁ��Cj��%8�`�d��-�r����(�1�4�.+�,���S?���%5�h�h��9�ƪ�W�y����oʚ��̡	X����:KXLٱ�;f�"�^�H�7q�|�6!��`8��q9C�|����n��Q-�mBEM��h�vtI��.ZC;���.��<d�j���l(���բ�Lv[�?���ޣ�I7Y���.�q�$oŭsy�
 ����Ĥ���������F�A��~4V "�]c��1&ѩ�
��L��;�,���0f�H�D�mN<j�:G��JD��[n�[���9�?E�����`Tb�:���F��閰�P=�g��q��ۚ��s����m a�[ۂ<��J�E�X[w�`�����+h�a��ti��p�� _�����d�������ZMh�����-��K���� ���ӛ�B�#1�v&��r5;oW���s��G&z���(�����w�+=
RB2@*$���"̷�+�����S�� �VA�y�tϔ����D��l��$Cf��p��Ғ �_'��OFr����5��r�!���:S�d,���u��u`s2F@:�� G!_�����v�☽�4�3������I9G����
w����ɂ�Pf}��fi�F��ḕ��/���T����V�[�f[JG�cz���<����,���mj�4��X�%K���2��x�hgs<�x�S�G�g-���k�^{$�z���&ئ.����J�i�[�~�4��C�h&��?V`�l�kdx�Jk��� 9�eЎ>
��N1[D1{݊��(���D�b�K�c�H���ǧ �b�19�fk��^4��"���������O�����H�ƌ�/UB�Q��Jo�-�����^�������zzf��M�_��Uj�����ᾖ���I��q�Y�ݯ�z�
AA�S,�jt�K�E�����a�h�i2U��!.���F�d	k��FM���ʾ�����A��w��]9K�sm�З�m���cQ�>�sV* ����?���1��a�:��O��	ea+q�-E?(�0���{�,4��e����V߉��do��H���{�}>)���u� ��'HU��������E�sCVrc�\E!���WE��8��٦�q���,�s���?� �Rm)��I̊n�g�a �'���e@�X�&���&�`�͘c��j�^5�o6{�>���;y�4$s����oӇ �!o�.z���&�(MN���~#�tqnЧ����Ic�����R><���п[F�gb�=Nn�[�Q��D��������Y4�����~��;RA�eZ$�//>�n�2�*�M/�@�)��qE�1r(�Q���G��ɈM\�����/�VN'<� g3Y`/��Yo�i
6��#q�t�K�x����/�3��pXdn��x����;v�{�vY����� ���!J.��wd�ۀ)�Bs2&tQ��'K=��(�*��M��Zao�S�z�<�X�D��O��s��L��GG�4�9����A����ؓfm��k)<H��7�m�6#����!��0L