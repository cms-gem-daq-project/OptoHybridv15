XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ĭ���"������ؖ�X�;��?x]e�o�]��9	y��q����&Pt�s$�s�Y��~�� �!��]���uh������p�e�ܰ�hp��9
d�j�t���_��ƌ�IDY\�<�F����kg��m-����yt�!Th��S��&̉S�ė*ϰ[��_�3�I$���38�񁥂�b��3)Cer�(��|if� ���0��Gno�-{�;��\��>��!�Р(3NlK��!�7-�7�Od�����$�GjC�a�!;�/���BS�'���amƷ2�Zr�\d�D~��P���ʭ��TnM�XGm�v}:9Zǅ�s����{#yK��18=P^]�| [�G?G�D��V
�H9�l��+G;��l�������ؗ\�O�l*�O�.�JU ��}<��{�[0x�3l�	F@${��$�~���,����"z����XGu~0��"G���@�0�X�ǅ�ؗ���;�\n-v�/ɰ��6���<ȕ *�����D�[
����hV�#�s�����*��ΐ�&@���u�}~k�W��'j�#C�h?5׊A�����<HJ��͹�.��Zu�̜g��7ҁN��`�i]�QQ�F!���8�s˭�1ћ�F�u��g��. 즯!�����*$�^*$v�Q�,*����b�]�O!��{60zJ�HlG�y!Р�f��Q�κ����S�O~M<�@�[J&|�'��tS	�%d����R;'����y~g�X>wn��H"�E_��XlxVHYEB    41c2     c40���G�b�}^���o �@��{H��]P٢��q���^�*��L4�(J����	@��x5Z�ͤ�k�6�#̑�^�57��e:ܗW֨�\�Pe�����;��"�/�k��o[��`�,�P۔���Z��R�@
�~'H�3�T�g��H]�M�!�mB� 9�m�] �:ߏΒ(��eD��V�sf|c�<�bpK�	3cT�\D01�qQ
c��Y���m��)���OG������m��A�ԓ���yҭ��+��L���={K�L�~(�S�ےie�1KTʸ>%�q��p�K����a��HR�-f,�8��Ň:�b �b�P���=��qP�������ny�A%chf��ۻf��D�;>\h��
�l��Wu���x��%����N$���ڤ�A���l"Y~2J)���.3,y�y��@��� �򏩸������<:o�������aj��XE� 5=�4gγ.�q[�7�Z����n�]Aۂ�3�x�̕��c}�4j����g�fq0�:�D�4E҄
����`�Ӭ\&�C�#Q��I
����|wB��;�gڼ�=�f��� �u���+|� `ԇn�/%i�z^�|�|=9�ݪ�W��*��"?��(�|'�xpܠm0����	���(a:��Ld;�x��:c~'��K<r�#���V�[S��<)1.B�E�^R�����({��Q_��jZq4��T��2�-F��L�;HEO ���^qx�$�a�K��&��L�cJ �c��2���8��o���A,�5$�h�p���i��\vj�1^O�:�x�SJ�1�?EvX�TE�	W��|:���UU[��u��(3y=�+\ة�Vb�@��f�S��������mFN����8&�s��M���ZEMæ>	�� �F���B8X�fw��FM��Hm��Dj�st�:�8�63D�])<�e��)�nɗ�}�{b�XG���=KhE�[���NX��.DG#@�Fu$q,'����l���������U ����Ԙ�L����o�� K@����>đ����C^i�[!��֠1}E��p�	���K���ݝv�]��<�o��b�MG�#`�;���|����y<���qLb��d���\3���O�YSЙQ"���P�2N64�/�,C"�I3�	�0%�r۬�@D������P�Rn���L��g'MN�`�7������y�5��v��]:q���r1�����4'��/9�:��q���ꣽ��{=�)�r+��8�c����\��c�jRJ��͙�:�F{�l[�/�pͨ�
ܘ�	��G���w��/� AG���9��Xs`7ϧh���?�;њ�o�S� �޸UXv���#�4!������^0�r�|=�@�c�<���Q��b�uD�M���&W�Le���[�h\�;>�G_��Z~{p7x�-ݎ��
�I���\aH�9��{�����{�}uu�u�����p�:p�8Ε��\�D˨���p���78��S�C«����]F���b֙K�t�/X�t���	ӒL;-Yb��䆾�]}���2�����"D|�~6�q�2��f���Ǒ~��	��]ݱ`[-�p�,h�R���jtʱd��#��SN�=���]�ڞe�����r�=0[f�K�CE�������3��T:7�r\��:훎�v9T�~F+B��Ͷ:KdBVnD��X@Z��>;� ;������Mp��`^���R��PB����`>9�0�q
��ԒZ��Ϥ�sϏHj���3C�]�E�BJMq��R{YȖ}Y��c�p= �jH�C2�5�|��0������m�_yga�(8~~�u➑�#f<����ߚt�Pn|g�1ž�݌�i_�e��o�Nݶ�IO��|�9E�U������J�Uzt0���~9͝�aY����I�Ú��7�SM�W��3<�:� ,<�Z�V��p_��&���L�rcby��r	!������P����P���O�$���
��~�Lo�/�?C$���D���}����13~ۓ�{y%��`�	do��:��o�FkcB9�MW�\�YYl�4�!<heIk�3�C�T�S����/[k8�jyc�	���~��Ǫ�+5)�ڰ���h��^��*���oNe�[}Q;�O��&ۗ���9�J3C�`#���dY/�+�z	Hے�*��J!�,�D��긮Az?��@'�^������ >�^��s�DZ�Q�W�
�Ԗ������%����|-��7B������]�D���C�� J���1\��f���fN��:5�����IB��`�Mfi�e����:\*�&n'���t��N�V�a L��ә����I����0��OB%ۜY%���Ϸ,7�ES�<TE�JB�Ipf��z9�d�z���_��,��u�������wBufԻ�"O��J�\��3����ϱt�L,����3ucjt�.��C�m�3��)^q���h��HW0�R��+����$��+�
<�Í��e۽Eܿ�Q���=3a{h&V4���F�b�Ա�Ig;8�^�\B��P}w�\��[�� �n�(3Ap(�Зud��T8lm)��V�'���*��\� ݮRQ4��a��;7`�S4n�t7�1���ru�:a���p[���1�JX�/���b�k�E4�IpB�hA�Ɓ���<$��'����ʴ?��#x�[��:�����V\O�q���'z'Vz�|�_��ŒۏX�Rfݘ��;�G��@cb�)O�W_2<aTq�C�f�F���ǱF�td�a��4��+� -�zDL�N��) %�vSt7��v+�v ��ֆ��a�Z����$wZ��Rΐ���iy�_��`?)|�a(�V��fV�a��T���t��kר����-�L�AYE(=�mA��{���:���CpT�&������%0�a�X1��21˽I�b������s�T��i��
~B߻�H��8�6՟���"�/g?o���G����?�������m
���m�Vҩp�@]mRF1�Vr'�er�5Z�R�&����j˱RX�H�H��s�