XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v��Z.��0W?��,&�oo���H�HQ_�MH �DM�~�_z�e1��JB[Ň��D��H�'����z��q�Կ���ɲ�ϓ�tS�m�6�c���I�avE��2hg,!-$nd����>'�y�I��ī	Či#i���_�iS�B��ۀkҪ�3��z�\�.ǝy�������<�N�&������/IT��뮶���"���|x��R��K�YL|��"�nI흍���&A��7.n%4�,P6\�o�;?v!��C�?����ݧl�^ |���V��r2Q
�Z�Ѩ�fo略qa��K�B�><X�v�/��n�U�����pH�x��i�m��_�k,��)m���W]��r�ڝ-"=]]4�m���ެ��1��,�-?��p���{\IL�7�3I,��b�E�<E�#���1y���R� �di�Y�ks��|�b�K��r��!T�+O�(��8�#��	m���ܧ�{q���ߕ�ayG b)'ՙ����0sg��e�=�I;K =��� �t��Ea���g�	��C�?�/>����7��r�=��椙چ���L�c��$���ō�#˨nS�Vz~VtR����-�H��
�['g�\��_�Z�\.�K�I�K�6���r& {6nV(�u��`@ڏ��o�L��c��]�66�Bc�I�t�
{���>2���ˡp )���4jTD�k��m����؂��FyW=�k��_uV�����H��|;�%@��ϼH��mXlxVHYEB     7d5     300Ё���L)V���{!0 ������7�f#L�3�M�`�,�îd5�KŎ��e��$h�x�Π�KY�B]�syQ��:��d��V�'���m'�|(%B�EP�$.\:]q�2�5vd�5�L������ pЛr�Dl��uƢ�p��;JYr~�B��F&��!�q�����:��]WITk��,g�i�M�R8���	@�&��S�U�%?�����z�
��@�9T��x"<�X����ٹ,ǁ�}?4�f���y$U�A�y�t�s�Fם�v��{O�4��'���&KX5l�3�1'����1-�e\l���++�9j��#��z���P�D�d�Q��Y�^�y<"�=�E7�*mL%��x:.J�8bR���*o�{�$U<�<�_�l@W�ԋ�����:�V9xr�w|!X귂
��J̬��a�<^�P&���:�ڳoE��Bs��[%˧��Z�,�̻�	���R�&��!G�� R.R��m�d�1ֱ�'q5Z�xiy���;�~��{G�q.�*��:ds<>���k��}9wZ�����̇E^9���O���("2�?�����BG�r�B��; s4	E��O�̔EW\�ƃb�� s���]	mi?��G�zE� ���b�Ih�;�eľ:���B����
�s4~���i{vl&���ܠF�gU��"��)�#_"��O�Gs`_�䰮�l ���Jr3�$^�Ft��Z�D��5#�I��su4��n2����