XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K��,�h�
�T�\��ii���������e-�Ndj�҃�]QD��n2��3LI�6R� �'&?�k�b��0�n������Y���IV�- �:n��k$�i�z�%�檽���[�ɞ$}��c�{�?������z.���p;�)����8��AQZcNit����'�5G >�$�im�2^�e$ئ �N�J�ywnx�M�� ��P��������<�/r+�ϪoAC���<��|a�a�^�h��u�|�q�Cf*{�ǟ��Ukd;3F��L��K5�7��޵a���Gȼ��H�43D6١�F��e�R�B%v a�׳
��_��d��م��[�+#�9�̝�#�1䢢�vs����{n
�y�
�јQlDuF0��|&2w>5~�վ����r�uTlMQ�>|��Κq��=I���Z��q�;@���Ec!�)��$������� <}Q�ڶ��B��۶�jedE�I�z��Gк�u�98�R�rjJ�7�O�EES���9]��Qv�L���>��,��q�G6��s;x�~|U��%)]7.�8��t�A^�F�߀�
�:$��Gl�B�s�!Jn��o�n���w��
�����r�	���U�U6d�B����[��2��W��`�LO~�Z�v��>�>lJ(�� }��c|�l��J/��xPa�'���Bm�"�S�\^g�䑢[����Kp��X��&�N��S��	��i��b�`�D��1��{ڌ�b�xo����,�5o�XlxVHYEB    a6c0    1b00>H������$��+�BvFW�nG
���t�B߭;�pР����oX*M#�s2�Z�;�;�I� �ӗ� ;��h�}�Pht�c[=dc^�D8Aߐ���1��^E�a
n���,fm�X�j���a�Wt��$(&8Cڵ��X���0��,{Q�`�>Ru��0`���Ʒ��([���k!3�/u�M� P������7�NXP�~�r����h���~!�w�uӑ$��")
�m���|y�0m?�W�������QA��^��b���OnϘ���'��5�0x,����D�SW<)a� O��#G0���(d��I�`OMOX�r� z�������УA�6\}�-w��U���D�*�n!�!�'�^��am�TGX)�xm�SK�em��d-}D�}�e>�Ǆ؀�\�C���f�tj}��MZ�!��	q�4�#x�[�����"�	A�O�R�ӴZ��
<���x��v���=������g�Z����0����tb�#ً�6ޖ��zň���竭'�(�.���_c���j�+����V��[��j?�l���tד��HZ�'5�I�2�����ԟck9,b��վ�����X-��J��Ål���/����*�L<S��_�j��'���x҆�KL)��%��:ōꉟ�{p��A$��$������K��aF]��S�
��?b�Vi��|�2����4���U���P�tw��=|��Vͤ�]�S�;HvF ����u�\Q�h��YG,"�x� *t|嬹�jށL�)������7����y�ct��m�>r�JgW������x09��$8��J�qkg��Y����tN���I����}J��W[����1�9�炂k4쩐j��%[���hL�%l!�	���N?�#m�/0�ź�o{��:[��ʗ�m�z� �����S;ޞ�N/ϟ\#�f�W��3*�
�=���[.6&Bb��o8>��xXvz4U��r!���$�
� !j�9]%��:�j�+v�ԞT5���'01��_�G�'L6a�z�1���������t�G�5� ��,���q�� TitiY�9��%l�'�*��H�.����G�/�.K�h��%W�j��R����j�r�eP��w����hݏS+{9 �'�$lu=���n&2.�2/)KHy�l ���3Jg`s��=�20�����][�W��k�#������V���M���F,Ǥ]X ��ȵS�Ŕ�U�Ițk�:��_�ú�����M��W`Rd1{�XY�/��U�1�=�k=�S�	�9���̽'��S%��5�@�W�fw�*�#�b�5�\y��7%��saj�MKս��q��V�nl��*n��.�Ql�Z�D£A-�ʨ��L&��[�Wӈaя�R�d���W@6~��|a�K���*d�h���_�Fw����;x �1o�\��P���_����͚JG������}u8��Ki�ln�5T��;�����-����[]�F��MrN���=�����{ҡ}C��N}(��y���o��3O�l�k��̒��e��d��(͗z�z6���
�,~���\�*/ʹ��_�!]��1p�` ��FI�	|�2uWW�V�+ŤyO8P�a�\N��T8?��q�h��A��)����o�k�1��bL�g�b�js�wS��+����5�y��0\���?7ۓi��=�E�%�(Zy�O[��읇��M�V�FM�\�8�I���=mG�SNK>{�K�ϗ]D��s��wu>r�2Xh�s�:�֮z15X�Łw#_;��Ŋ/��v����U�����F�-�c���|~R�r�2�+��;H0xc Z�tWb�^F����V�Ę3�I�B�3d?��rD��8���OE�F��3¤����A6�,l �'�F �UMD`��|�!%D񱫚���g�W��J��S}J�ZgVħG���l��['%�bRì<����G�#85��in�)!Խ����C�h<l�_�?�E�>r;��#�ݠg�a����ֽD�0�����,���ve
Ok�0Uon�r(��mγ�� +�W=�޺�'��
� ԝ?��M��{��4���Yp$!S���Qo`FX�P��7���u=.�;e���N�>
o���J��/!�S�g�����Sb*�� ݱ���S�g����D���>B;1���3"� �*�oAka��M�EY��x�6D^�·S��A0&���]}�Z���M	�����:��n��YFՏhՑhS�?�M��z(1(N�����;t�6辐��k��g(q�N���3��F��� A���hs.��G0!nw��,v%1��Z*��`)�<4b��#�KR��j%ҐO�3���	�(�uL���M��+�ra��0�1��zϋ#�p��es�!�W�I���Aw�=��B��Ib��߱�ԧc\r��"Hm�b3'��������p�8ج'���
�����X���/9�%W:�h�s>j��4L+�������?> �@��{����{�����Id �_�ř������h���/u�����tj�`�� VM'��#b�,�G#@��\�}�8�0�]�fJ� i�<L���f�i/&�R���G����T(xi�u���q��{i�f���O�+}�a��P�a(B�b����c�����v��8�M~����F���oϹWV�"�d`��S�e�u�	�� g�P=�R�5�ת�ȣ�>�|'����C��󲂪P�B�!|��w+q�Ć���WFM�i�|�v�D/)��A��b��UE*�K$r����-�9���9�5\K��F���:�yL���O%���첰o<�JYL��p����,
�9�38����*V��R��G�k��Ko�m�T�զ9}�^���X&&yF�~��5���Q9��P+|��\��q*k�::W>���fV�0m*A!�gdi�+�MҺ�._P��(D����"rp��M4����&a>���:�����h!��Z����
��}�%�8!��N�ǩ|��N��@W}Ǹf�+� CI����nܴ���=TfP ���"�!UDZ?�?u$��1�x��UJ�}�~z��0"]��zS�
���N���޳�D���@8H�:����h`XPl��gOEF��/�fH���*×��E�/t`� b�i�tg篷�{�2�_�T�%�I�`�&=�*Z������1sGYܳ�\5t���e�DK�2�r"�y���l��/�=�Ͼ�$4����bx�B�3��fI%��ێa|i�ޏ(W9������'���P�,��:e�\�
��rd"n��-�*���X�%��e|%g�+����ߑ,�=W.Y��~��
l��ȕ��B�k�<`续4H�6���64�f�e����m�1'�����"�4O�R��3�%2Jb	�[�*�1���ж.��
<;f�ǰ��1ä�nV�S1ݽ4r���7�0�e%�:]̕�����ʆȦhY��z�Q���
�<�"�WP�r.�b��az�G�Yx��:�6?i1�����9�g]����p���z�`����Ϥ�%��I����B�y��_`Z�����0�U-��ۤ;��dzR�oBj�S��ri;��3�Ii�e6cN��ӱ�8��	�io'�A�/�\��S59<����T��.Pu�W�-�>����}j<ґ���S���7����Lv/�H9����F��r�Lo<(�o ���!Mp��K��IL��0�ts���%o)��ҔIg'H��������첽�������/��`E��^��K�y�+u�u�S�۪�PgL��
��o�����hZ=A6	9�;@��2���׭_�э�Y��|�C�S������TXں�3�9�6s��&;���Ͳ�S#'�+X'î�,����F�?]	M�댘��_�|G�Cur2��88�F&�K���F�]���ݬ�r8����i	��g�$�v�f� It�g����=$�cn�)�<�r�!9Ԝ���bR�Y�'��e��4՛X4���h8���&#�6} ������������>����1�{�M���hrVVlޮ�t<�2uri[k��0��YA"Ti�[K֦�E��Ⱥ�ӷ�`w�:�Ja�\nz�d@3g�K6��O���N��!QV1�|���1a5m�e��=��>��⪰�T���?�tN�_.6e��k����xVMd�y����;�U����IM�3K�Υ}�d� vf;A��;�^�s$$R>y��(�3.�8&H�:B��R^�A��N�$��+�/��b�Tb|��i~K��(c�U�{�\|M<2)W�L�A�3����ɗ�t��M�k���G��諃�t�y-�˫A`�+1�\m������zh? ��*�=�J���
,��Y^��4��� �.༓Fdt)B�����cX��O�ZݨE[��K�������#RT�AY.���\2E�rt�jx�,�t���1n�*~�4��۬�����{ݙ
o��Y�@U6F�m0���q
�=�?���?��]��������@����$�����(�
���Un.�ą�.wB�%@m� j���<,�<�P|/�b�S��~���m����#���
D����Ș�B�q���oƣ����~.�j��Ȉ��X�.�/���o��g�ȗ��t/c6FA/�a���M>Ѝ����nE[�|�(�/��z��� �袎4���N�Qz�E���3K�=ˠ���ՊɈ�pka��s�������ņ�E7��Z����?��m���76
W�_`�媧�;����;����{�,���R�O��Ī��������q�����y	���j�*W:�E+�%]e~$��������K������?v,��L�f%���Л���.)��Y�t��(ūb�w�1�OcЂ�|4 �����tZG*�|[�l ^�Ѻ�ԶP6,�r�� �f���rU���p<���"�tpWʲ��E�hS%�SN8P6�@��������?ڟ+י��f��';�A$i\OM;��^=[s�	���~ڶ�~�e����� P�qs�Bx�FWa�Y0w���&U�
����v��j(�TA+B�̀�خS]*$���7�\fқj��l��,��j�������Q����y�^A�5�&�s�]q;0k�z����0�$�,�I1��:���dE�7�:X:���J���,lj�֨���[5��OOg��x=���^��s��gn�R�
Ǐs6E��@�~ȱ��V ^��zm���:���[��1�,����`���"A߫B�s�_+�s�/z�j�1��a%�XMpU���/	(aN��vwơ����OL��Q[�=�/N#��Ҧt/�c�RYC#�K;[]F]�j���գ|���k�)��u[i�
�΄S�ச�����4���Б���-wCM����<�!����� �#�l���]�݁$0(Y���s�xM�$�ֆ՗dJ3��-�����&w� �q�T��,��3fV�9!�|'�!^�kǠ�2|�v8q$��jӢ�d-Jk��=e\��ȅa0�%�����B��z�=�S�}�<��<=7ER���!n�*��ꝫ��ۣ\���ZM?:��7mA_}~�l���OG	t\�^�r�"4	n��6��l��s�=z�$L����@��e�k�����#:�zVм�nV6�Q�H����#�Q:5h�+"��hE���=��h�BF���3ǖ��_59ʘv}!���3 h�[�KHt�9�[��B���Z�s���@ƫ����b�\s��m���ñq;!������B�Ľ�K4M#e����A4��p~��!����/��^���_-\~F�[7�Pz�%�� #�ڨ�@���<Q�B	L'1���@:ũ�[�H\ܗI��;_ʄ/P9Ͳ.3
���Ga`����k��i����{;��.=l A,ǆa8vHLS��")�.d��:i���E�Q�܌<�I�wt; �A�C�����u�`�����d��K=4�� �2�;s��UNe�W1��d����~��߼͋�@
i�����W���ޔP¤�R�?n/@�z��}=������i�k�u��DWl"|�nT��,C�-���y�1�S�d�� d\��لT"sx��N�r�\5�͔��]F���T��!������*R2@y(�Ϩ�$0x��~x�Z�0��WM���`x��b�nW���:NKs��.�"��-�ȒL�q	H�Z6�̈�Pb;�pa�{�C~s��z�LV�jUV�3�,h�yH��Ǚ�K���E*Sp��[���*w5��K!�,��^c�J�xa�25���*��\w�3���^� �aƟ2�@���X��^Z��_�me[�7
S\�8��_0���M�g��:�QL��΋!�8BB�)s/q�.=�� �J��<�}�)u{���[G�^$��h-�ˈn��M��%��"ͺ�@k@�ȑ#��!���y�Yç{=]m���|GP�1�T�Z΋6��73���o�I��}V�0������%֒��X��yx����2���!
���R��,���J>���A8���$LO5 Y���E��G'���xwD��b,�#$\�v'I�L��,�oRχ�|k ��j��n;��bT�PQ��X5�(Ne��le� ��|��߲�HCvi��G��Ŋ�aP���#�P-��ʰ��18��P\�b/���Qg&�X\U&\�!j%]�g?��:�ߺSd͟��#��M�