XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����H?h�>?*:*_�#��%��"�Ş�8�Z"���rж��P�Y���p}�bXv�~�/�t@M���.8k�$$��É��%`�������F�y>(�_�펧2j��wЊ��\��'��uZ��LY��YOR,E��2s�1W���ČM*�p��n �6�瀨�~��@�6҆F������.`+�CS��G��2{s,����q����B%���@��a�\f���}� \N�̌	��92{�5S�"6NǇJ(o���T�Dxk@'�>��%���*���&����'��N��G�DI�*�_�Ayq�W&�Z��rw�s���1HU���gM�"�v/��"m/b25�iI�h-��j�6B+s��wQ��ɘ��w��G��v��R�^W3��Q'�y�S�����;՗`����,䷕<sV��@4�?C��L�N�<�4��~%�	�P�G�"[/h��U,�-?���I�5�l�c�A�3��0���f�{� ���:cΧ�1�'@����Lb"��I�&u.QO����[U��t�y�_+�o���/�χD��8�!�׀��beQ ��g�<�.{�Bj�/.���}E.0�Y��I��`ZRO V�"^�3�di��\@�dH�"}�U�rAiH��M z��y���_�<q���Skw��M�G0�eWOSM��+�Q1�Y38D�5*]?��^���9\��3���!���U�Tp�e�׻_g�qQSF�2����|�̳��8q{��kfC��W*XlxVHYEB    15c3     780�H�%N�S�)h�l�������aU�bA�I��D�[ח[�l�$��;��"�m�ʀ��G<C&!�[Mb�\ۅ����X��D�2���Ew��G�b?�%I4�J�a��IX~P��v�?c���1Ĭ�!�=0��C���x�������w�%�-"��ȴd8����u�D���C�n�;|1��N��*���$�j�!���Al�5�ԎP��ω
+M�R� t�%N�m�x�sI���D��J��T!�r�6h��*R=3!�~CU6�^[�]}�IV~N�Oӫ�KpP�7f@a� �mK��D#)�'����-$�MU���/b�P��H��^(��- #��NǦ�L��XF8L��~s_�+��ؙh3\����îޢzB�3�֏���5R�E�3��X�gc��Q!�IFxNR�
	��*
�������Ĉ��֘&F�g�U`��P��B��[��2�a���)PՔ�j������3����x#u�mr )�ǘ]��L ��}���ǳ��Y˂i�4�&�dE�G� �l��P{,ۖ�^ �6�]}H�`*|�Y9��kh�OD���R<��5f�S]ej��e�x��x����Q*�FH�?`�ޡi\�Z��2���Ӈ����ԝ������?��rc���;[�C���m�
g%*ʁ��:^�0a�H��ҘM��i��PP�;�Z7�IRV�,�*��f��u��_^�+���=�9��!��tl�#��W ��9��P��o��뀐�/A�|�G �V�v9�b(1H&�Գ��<2�\
�$/�"��K�tZ�$�����=C��
xѵ��V��()�,�7�W�3.��1���(K�wFs��鏨�]F>��bv ���!��ڍ�.t(��_j���5����Dq�7�@����
�]���O~H�3yI��R�g�N�8j�/�
����+��]��r�ps��[ֻ��̊�7Ŏ��F|��I�*��Q��x��6�1�����ď�h�\j���l�&�W���Ms�읗�6o4�K=�$�B8�6�]-z�ښ��9+˶Y�����G0�ֻ���^�}߱�(���-x�Y���WA ��be,i�\9 ������G�4.��yZ����G$�I���BKѮ�w�@�;�ϔȱ
\���?�0m���r���	�MC���W{���Ha���gb6��Զ3�tE��D�i+ۿ�N�V����7fS��\����W���n s��U⑴���Q�v-�)��;Ug�@� x�oS�*7�ٕ�0ՙݍW��ŗ��[�<4O�����1&4.E�
��lI�D006>(9l.9O\�>}v��?uo��P�N����րq�%��xbK��!�fl�>�4�^�8���E�E�Z9�H�7��\4E�-<�,�G�~��� �>.#v\$8��}\�iF{S�y��{c޷�ߖ�&.��l$S0@J0���F�)\Qf�*����y��YgZ��H#~���'���ĵ����O����J�����OM��E�H��c;�ķ�d�(�8��#]9��	C!:[5�{��vo ӑ���s��DiB51I#��Jz9�����!��6	��oh7iY�v�.��f��0�Wh��3�F��Sy'�/�(��2���j�pU:��19<'�b��YN9���Z?1u�������<����]������<����7��F:>��*X6�Lh3afi���4ۑ��c�pi�ԇ_����d��p��Y�]_���!1�=��_�Ԅ�S<@I�s�6M�kT�fd.���N�B�~���hl��7�+�R����X��d�����`�/��b�T���0��z� iU������8.1),�M�S���w֊¹�W"�,���3�X��f`����F��1�+��z�h�[~��	�daY�