XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ӖL��	�c���Y'	7�zu�%�Ol���'���Ձd�%�
w[8����0��r~���������󡆡�s{�y\�%o+-a��e4Tf�0,g�!\�,�X�D���mb�jNk��C��/�;����/�{�yĦ�~3�W�ܱ� ����>�b���t'i\9����I��_���|�r}��� �Ƭ*P�avfQ�1]��6]��;絭�_Ō�qj�'�v�+����Nx̝����~��:�9̊���x�oz-�S��2깉�l� �%x���JC�*�V��c פ�6l��7��!���A�	8��A��T�XvY�+p���a�����`t�F ����}��%\m)�3�����>"3MP��aSj�W<���m]/L]����p(a���ݒ�c��w+]ǳ�6{i8�	
`�*p�?��Yr�?!H��R"����8:PEri�Ӹ�$�q���t,���4�j�J����۵�_�R
~����z�q�?���{.{�J[����*S!?+�+�V[uE��P�k{J;��" T�JUZ0f%���@7��t�r ��K��o
���z�;���q�a�# ���'�l,���tf���Y\$�� Ifx'@��AeQ��1_34���8\\?@.�T,�W `����,<�AW�{D>����!RR��a��,�vЀQ����ZV�w/�5̎2�~��;�I">�\���U�=��	��C�F��5����v~�����q�7��u��/�p�bB˶4��&m��xE��H2�XlxVHYEB    2d5f     800r��<�{��b�s�r�+ˬڢ�mDV�Z��R��%?/xq��q̏M3J�s[�΋%�_�AN7��>f/g[��N�ױw ����5������B0S,��d�Yc��K��cf)�<(v�u�GpIV��S�HSq(��{�<�W$4h̖[F�A0N����	���#N���ٻ�*OA5�c-� ��[`C�:�S���@a�/H㹯�R�]��Q&���0G/���\G����E&�A-s�O�� ���
�R�z�jQ6w��M�ø�K8O�4D�����@���, ħ�@$�ȘjEu����%��9Fs�;��REA�sR*�=��1���k^L?��S:�����k���i�3�xa��)Գ��f�b��p��²��1�]7'�u��t��W��y����XmW3�K"����Y���1κiɌtYN�H���=+.~��x��
��������Zc�����d�k�F{��U#�8~�j��:��m1���{7��<*�smo�n~O��n��B��B�%��|��h��q����a/
V�4���l���G��f��v�6I��plb6��?�aPͼ��l�5�A��s�d�1��j edt�I�]C���f�K�}֬�l�
��Ju*�T��s�A�`��HM���sÌv��W�̥�J����jl�B������T5�,3���z:a�	{��a������э_J/>ģ�M(��3�B���(�d�]��`<z�?�'����PN�n�:G��Rj5RUb�x�Vb�Lc;�еe��
�z�^��FXZ�[��OO�;m��m&��8�I�7�.U�G(:╫��'p^������3�&H��Y%������J��OQ\��R��S��L<4v���t�Li���>��q�H���	�E��!3z6y�'�+�m�+6^}͵m	�4�NQ`ӯ�;���l�����WP�]�#"��>I,��Ƒ��R�r8;r�~w��8�2���+�׌���i�k������%ڦ��ג73?U��GKj#��ɸ�O]�aƪ�*s̸��}��`Z��`M����������>r��x���]��5��/��"s)n_���U=��G��A���wf{Cr��<����b�lҮ��d��	Yd�1j1���,������S+2H_x�f�q��Ma)�5�ý���ǀEvoݠo�?VFv�s�cUm�� *#h�yy�U�������cD��:	@.�	1(Q+�/�̶�(��(B��xŽ�	���=l�@��`-�O&��m������sU�SY����#�sq��C�A5d���C!��)kˊ��2��i��-W�s"�e�l�v��Vc�/��6����8=CU�Eŝ�$�����X5��n�@����a�H�o��<�SC�"	Uݾ|��I�Bu�K�3�p���y?�Rk0���������W<�s_�0���b��d�@�<9�ز�'�O�IȰ,3����}��PŚ�?�&URu��H����cP~͂7��yj��I�e8�Y��:����F�c����'�$f�`iO���b�]��!V$Ƹ-�z@��eB͗�x�1�pxي�l硥�O�B-����'�"��{��Z��GD�a	ؓ3A�Y�X�u���
���]i,���~O\��`�� �� ��qD3vX�LΈ^j�?Əj�Q�5�����Y��)���
_�J>*�7[��?$=ZK��Yh����~N���at�պĎ�N^v�r�1.���BT�2���������ܝ0N�8c%���;��r��.CsH<�Ƃ\��'���9��ʝʇ��TC�ª�n���S%`֋,y~"�Ч�M�d�OF����.CQ56�'5�"(I�t�jc4��v��^������wZ�M΁�0���RUd9{������dfN��J%�N=��~2���ŧuP�|\��W���!�"��X�"<�fG�'�	��E�w��˫e����� 73�