XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/ʛm���i??��]Z�>�^��(c���v�o�>�>@r�a��/"�b�:�VzfmO�� ��������/�J����9��ri;�c2����
G,�g?�3u�'�f�r�;��c�-Q�g�p�O°(�7�$ֻC@�X�i�Q'`)��M����2�(*�ʑ�R�^�!ķ���l99U?/!6� w���������%ꁷe��,�5k�o�l�^P�V@'���9�'���ۺh"�������>��7��H��<�Z�ЂR�9W�v�5�8ʹ�&�F���u0U��hA��<�n�H���Vz�e=~�5�u'�-w��xLps�OT.���)M@��wm]�����,��� jj������E�i�����<�`�j��[gmW��3L�u��IE���<���,\�e�(��H�գ(��Ĉ�(���呇>��	��bF	(.����m�{���\��nx�qq��S`r�?��>0LE���!�9EL�5NL׼��gV0q}�&���N���2���F��Eݪ|�u*�w��uA��Xn	�"�'pι|�{�m�}F/�34n��dh��r�;��P:������'%7{�Gg(7�N�k5��.��S@�T�[4�,��p�jQ�P�����g2�KH���(R�N �'��f\Z���u�пɁ�"�{n����\��M��F�%֘�eK=M�"������Wx��Q4m߼���gt�M�#�ٰ㔽���Z�'���q?ޜX��`����]nXlxVHYEB    6fd8     c30�=��0�Kc��@�Eܨ�<��'�9�=��K'�˛���ij�vxi[���l�&&e��r��R9-����z�f}b��tJ%���������<R�l�G���곌��ئ�߽��IJ^!��~Σ9��9_'Lh��X!|n�Y������x�g�������u�%��:��D���P(��:��2*��c�(l��jO�c���s��|�J�4۪��B��!�{U�ұ@�MMj����"��B�L{�h�n2���CP@��V	8��O��]Xa(�HD��E�`�����Bq���5���pje�`�/�����YZf��'� (`�~y�EҔaoU���yy�S�a~>+���?ը����9��=����sn󬵣+�ϛcɢ�KZa�윎�"�P�=K���~F��'�����"w�#+錦,��	x����(�U��BX �}PkGt;?Ś��w��OU����n�.<o�R���A���6�?n#���e3]�l�B��Gg.R�F qqz~ ?����<�)�@9%o� ���=�'h@�s[*zJ��z�<�ֵ�A\����61�0¡NKG�]A�~�L�kʍݙ*��xC,�ٷ*r{V섟: ^�M뉜ZRc^��y,�iA�(�l�P�o3!3N��F��f�K�XO��� S3�S�Q�H�7�ݡ�o�80�ν�P��C�ɪ
�@\�t���_ò�m������'�>��[�{A���Psa���ࡿ���ϯ	 �}D!#�	g߱W������8�m
r��7�̒	B���H�2{�7+�4]|��S�!����hQ�i4�䃥��vC��GcY��N��7G���a����]���Es�E��G�)��@`����j��7�����%F�v�8%�+6���T�:e�s��`�(z2��b_a��(�,�f�]�>�WRк?L+hp����UE��Q�,�௏�|��Z�x��f϶���.D��aKI�P`��&�%�=L�%%4x�貶ju��Ӡj��Ys�x��g�^�ɲ�Ǭ��U���`_c��Q F���T���Zh/y�GMq���7����'���|Xt��p�1�l��3�
~�\�����@g�H=Dc�}���J�^��N�~�q�B�4��n��X����G ���ɨR����#��4�G�K���ޜ����fѪx�C$��x�C�];1t��Ϗ#R�Ҡ��n���j�l͸$/�3���h�������E��	0ihi��#0�_C��k<*�ҊdqK�+�"�\���x�e:����� �6�ʲ��˜�Z؎d��[��=si��muRO����'@��M��u�9����8�H�*�F�(*�}Z�|�H@��^.�NX�SDgj�`�T���Oa�y;Q��0�;��E�#�6�	e͕�n ��=و�s �t����>C��>G�?r�p�@ٙ�C������\�iAA��t�	��������z
("v�&���Գ8�b�ڻ��4r:��Ü��(\���0EPM�yP�|l�!���bRW�$Z|]�Ͷx�K��)*"���U{��)��͍�-hQi�ka�s����PQ�9�G[Ҍg���Sqb>p�O���=�Bɯ��u?�Y�efi۳	���޷�Z�[_2��;��f���]^f]�m��}Z{P���5!�$<��bZ��ً�֤$���J���^�o�l*����æ���{������f����g�d��5G��e�
(Cg�j/�\ja��.�@Ģ�B�����fޅV ָPH���,#��e}���/���s�j�*�5p�cYXB��^�ݶ�@�C�Ĉ�B�]a���T��L4���T%��3,�l�Z��5@s\����_Q�t?o�/���#}�j(�����]��	����n���Μ @���1���V.-�S?�d��0���M���m�Ua�+T��4��9�����9�o\�Y  ��7(��1�
&GGT'�:�>���	��{���y�
K1���I����	&�ͼ(�s��wN�5��N$�L������AL\��X]����
1�����+��N��2vN}��,u�e�W�m�L��U���+� �Y(Ɍ�N�c$���g�|V� �S M�(��F�$u���u��0�����?ˁ��KL9�b��Z~�<p��݊��3��Ji��3��q��"���i͵�#��h��q		9n;p���y:�J�Y�xx%	��f ���E����:����V����y�f�5���Y��P���1d�~P���N"j�1����)3�lR�#n�|��4��KO\�<Ü���(-2_J=�����]�v����a���BFV#���p}C��j�]Ҋ�Dյb�$�ЀR�/��3('j��C�u�/���p�D�F�Z��Ӵ�TrCV�8�l�T�&/z�|����G0�lz�1޶#wLN��981�Wz�/9�t��,��/K��?�?3�{83�.$��� �=�a���B��0�fs�\;ʉR�2E$�U�#hD/- ��9��Dd�z�㒌c�.z���}�-�[���Sw�Ͱ��9o`�Ƃ��C85֕�?�/������m�᧡@(�@ԧ��"���;�4woIi������:r��0��#���I��h�}(.����p-��@�qz�u��_�la�y�q��	�����4�~9ܽ@
#�,)i�-/$�ݨ��6!~���C����җ�����&i�'�,����6<o)�J���\�\�a�ޔK
�k��XyP-L'�6T����mb?�� w�ɏ�8Bq��]z�M/�� k�|=b�Q��/c���a�7�y�!V	`��f���>�Ҹ'��݄6�{��Irg ��xyc>�>3 k�Ouǅ?C��7ݏ�z-*�Ѯmt"�A�q�d$��ޝ|/���ԅ~CV`ɘT�8�	u������u����!2+n���X�q��&,8���	f���s �D@짤G�}����P�JDnN��,��h��!��׸:��T�ܿ�Ļ^sc?��Mi�K�26}ļ�5�2Cl