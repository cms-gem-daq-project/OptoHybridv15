XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$|
�G�3*�{& �'>PI�UUÊ�8H ����� :e��{�b�\��#���y*
��"�ط<���%RW��SUz��qٟ	,���,a ��޹1m�s)5���AԮ�1y�d4\^���^(t�|�OT�F��[�.	���"��M'�e�C���Rm��}8����F}��?�0�J8~��m���9y�)cl����.���)Dg��FM�����<����C�t�R�o:/�	<����g�.�H+}Gjs�+!��֛�b�.�ؽ䧽0�a.�I���2�[��*Ɂ'�p��{�kWf�P��_�c�F��9���L���)���"��.����ȶ`�� �����0V;�*��J�p�i�D�gC�������余��XdRZ����K��?�}���Fh.�����Iy��{ޝ���;�̴	1ܷp�e�M_Ӡ@���F�e
#Bs�oS\Gg������y�4�F��{�C���Oʅ*��Z�f��lc��Ǭ]@�;,2�d���O�Ҁ��3����k{X�H�û�7�s�;l7��E;|�vL{m^�O{*��9�)�t�ݩ��]F�!b��8��L=R����B��P�����4��=Z���u�O%R۾X�����B�D�m=�6�ێM�S��;XC�kB\��Q�⥆�8k�����
�;�oDN�ޒ��dm�'�!2��f�ҟЏH���	r��"�����RQa���֑/�|b�T��hm���b�+��!��O/�$�� Qd�iTXlxVHYEB    78d3     da0���,������gC�)�:�Rhم�{�)��:�XԐIjoi��y��� xsM�K$��I��r��a�J��������)���U̪3�s����h�d�&���z��\A��s�&���/��o5�M���q��,14���G�<��u��,�ة�S�><��#���}��x-��*��?z+��HoE�|9I>�L�4���/�-[rt���"ߥ�mt��L\���` �D�w�e�b��8&	����ORA	sK+���M��NC������q�+��m�]C.5���(*�O��t�r���_S%GP�w���\p���#�l�A������H�`���+�'IzP�@7v�"����0��L,ʼ���9]___jߡ��$L.
i����z]e�'�$\>d�'.P/�8� V���	�W�8;>Ѿ����-�Y��71%6�<�D�R�+�`&l �;��"���������|p�:9Q���V&��&�kZxd��ht�!�d"�� �T4��3�֮��k4�r(,�fA5���$hϏ���9�F�Dܣ�Y`�3��#��%�ǚG$-n�������Ei�(�D�?y)��ޔ�O��F/�����P�J��2�	U]W�魳�����},��z�_N./:�A%W���F�8��&�\�nj�:�S��P�{�2�7�b��u��0W���vc}�i|���1��_w���c�(��i�;H�58[?�9H�
9�ސ�k�D��&���Rn��Xk�DA^�í�4��~�$ya�i]1sS&5�nP���ɒs����.A�]H�{�>��u�r���7�fK=��DQ��<��fM���9��\��ԽN��A��⾙h�MBx7��������$��u=�p߬&����``�� ܺcs]���葕��pl١{�><{N(Ժ�W�[U�UXP���,��-I�{�8�Jd�!k<�nV�a��څ�=llQ��/o��3R��-3�-Oݼ���>��Ƿ���+Y�k���ز���mإ{XCAE�\ ������[�gu	"��q}t�b�E<.1D#�!��룾&s�Г�6�@6Gi��߱z��*��pU�x���y��!xnI\��sFʯGb8���eؘ�Qs����=Į��X�3�Y�-�e8W��򰡨!���H�G��n��
�g�_�no�hiC�jYy0P�\2�m�\�����}�߃W[m�ΌЙ�w��<eqn;��%3gϫ�ո�<����n�gS�r���~�h�بx
���k�T�Ѓv.z�k�$�48RIX)Ak.:��"��v���2n���ߵr�$�������I|民G�בR�)'�m����y��p�x��5�~��U���gcB���$g��Q�(����^1Xt���
��:�k��Jk�^h�U5o�5E[�!&݄� oF��y��x��\�,s�1�?��:Ρ����>�0-���)����Y���K��31���!�2���x}��n���F.�{kP>�y��,����s��F�;5�'��O�L׮hjnE�P��$4_���@��)"A�ǼIy�#�|Ih<�&G�c�E=r��X����-��Bu�573������?y
�J�K��;EW(���\�G@�X�mVׁo 2��X8��o���~���ml�&ڳ���U���tce�J,�d�-<�<����x�gZ�ȣ����N^Z�J*_i�-���a�9�U�]��w�X��]���WJ�F"D�Xl���<�)��:*5�UK��@�Y����T��>�=wB��K�{?�Hyx������y��pF��9,4�oe(!<B��(����|�������v
L�������o��J��%ϭi87-���JU&98e4UBHX���˵&�2�~��>cz� JG����8&�L-I����xm���<-ZT(�yI�)�?�b�_JuD�@�ʨD8��/�@rgԤ��Ϟ��0��n���d���Ff�����}� ���q/>���	l�-��e�1>������0��҄�N���9P�����k� �D��g�`�����`��C�f���q��ݶ�s#G�c)�~�n;}���H<�,�Z�-�Cg�R%�8��"���'�̄��8��^����{ZUA%	w�}�
-^�����+��g�iC�5s��4����L������ę�Gr�sV`Վ��Hʁ�U���P��MS����6��[�(8k�N7����.LD�Xޠ���r����G?^��"�S�rb �>�ۍR:�=�П�ݕ�1ow��K2�&����	1xo^��]�,��q���>�eHD�rW�X !F��|1������m�B���`f�K�|�y�%\���8�B�=�Ux�5�	�8�_a��:n�m�\J�./3��/��\�(��ufn�?q���v�(��w���&����E���>��`^��U��z��Ik��GT�<��+�4�[k�#�&�n��9:�p��°��e��t��f�ozC����j O���hd:���6��
w؁6�׽����x[I|�	ˠ�*�$��Gǒ)����V�~�%�IUr���4���h�.t"G�:�\���dV�]��P0�7�^(�)\�E�k������Ey�ܠ5Y��8����0�	O�j���~;."H��1�GFٺ�Vd%�GX���b:�	����e��`%��T8d�����n"�4����;-��|'�Y�*�A|�6~��I@��R��F��������á��@�p�2`!�� ��VM+T	�?g���]X���6��wF�3�xM������m̩�q�ҋ�HB���Sƻܹ���<E����-�j�&n"1;."����Sdl�_h�v7��6����uB��:~�o}�q"#�&���4�(QB�>�)�;��������K�¨a���ts����Wd��!V�RZ9h�%�m��l;���R�{��~	6�Bo��lMi��{�G���x;a�������?@]��u�vQ�PT�{�S��kGab��s�o���ú܃&�\��<De^�F�����#FߕM��Xv�����W���W )fr���ș楫��Z�p��ӃQ� _��W��*�Ua�5�dKg��d�-!Y�����\PT#�	�=
���N}�M?՝��W������;rГ�)�uC҃+�9-���˳��?����С
��Y����0�<O��oE@�{�JF�}�0r�z
@�m�޽��ߊ<�- ����[3�("�
�\ej����I$�}��l	�g��1*W�;|_/2���2'YGr�rY���.�VfSXp�:E�IJ���]ohLk)`�z����_��bPq��#J�t�b��\��ɯ��rV�Q?F�"m���h�x&_���]>��O�x�=������y뜵
