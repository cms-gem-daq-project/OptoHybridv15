XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��%�.9��o%g���ЇlP�\m�ԅ�+�_��h?ܙw�kN{|�P=Zy7�ne-V%�<V�=Tݎ�?�d�Ě�j�E�U����x4����Z�r�9��u�(�ڈ��	�	-��mعw�<��`٘ڠ�3�6�Γ�
>�䔯��&M��Й���Z}4>����\������4(��@l�7٩,�tK0��x���;�W�D�Y5:*7B?���\#!ov��;�����4��S����4G@�]�s<�;_�t	zɽ0����ܧ�W�j��4	�7x(cR�Q��M�}��
�~�	�剦�����K�O2{��xd�Y�_��J�kɄ�����E��V�i��@��q�����U�s eԞ!�|Y��s��5T���R��	tg���U�c=
�+|{;	~�Ș�ZJD�%`p7�Sb+�hf��b�Uj+��I��v/�^��D�"�D(���5&Z����=Z��6<� �pD��&��>}{0N�sL猷ɠ�M��<���C�w���$C��M���G��7k`�휚{{}�
���A�����"� ;=�����W���Xm�CxN�.7Jl��ə=�֖?uV�����R�r�Q��{��I诌8K���K'Ϯ�nﴩ�AO�w����� ���3��J�����B��9�}˯L�aj�pA:��k���Z@n� K;�Ͱ{9u"7����w�@8�ǔx:-{��eto����/��&����s������dt��/�;(2E�'� $܆XlxVHYEB    3a1b     d40�Qt��ϟ���B��-O�2d�N�x&}���q��r8��Ji̩:2i�Ō�&R D3,�nU�T����K��۸}Q��u���}@A�E�b��Ȳ�Z��sj���r��j$9�/_ /���q=�l0t��|�ّ5%��v�m��R�UrcU�x�^�ʿn�]�/o��fws����J�Э�U������/>.�:��.� [� ǯ�sxw���#�����j�v�T�hRY��f�-I ������LK�C��j��C��Z�C*

��Eb�WDz|A5+?;@�����(��`\�؉eI�|�����5����E�4nh���
��Lk��gEO$��4��\	�"}:���
�J��ǁ�Lk���|�ݵ�v�ً���]���A�y;\ԧ#�H�B�YE���
<���&V��p��es{-г-y�_�����ki�a�B����#R��!*��(��l���k�-`t{�������ӒKy�Ԛ�N�5^�e�B�.�sK��ԧ ��9Ο(�h3�9�� W�s�Nt�$�,dOv�Er�B�R����]���8�vkBcc��*��'����L���{5��������s�W���`��C�j���q	�Q�G����W�
L@�Y2�<uY^I�{_�b��
�u�	�A~�GZ��&~.�1ph�]0�*����Gh^���
��0�C�Y$�pRG0ؒ��׈��;��\舋�QTjJt���s�W�X�Hv/#qC�b1%U�"q��^�6ߤ(��Bg4:l�SW~2O������7�?׮�wY%����ڽL�5X"b��W+ZiA���[�CL�A��u<�������̧3�r����T!���w�-[�6Ao<M7yT�$;m�B��a�4J��&RTT43�y�]-�Ch� �4ϕaR����@wC@��$#���";�rVIN�~���*�}�S�:��L�0e�<��$�g�owe�W�i�V�w������um6��FB[ٮ��ۜd��#Qa�#�5�pQ^Aiת��[6TcuEx�T���\�ѩp�s��[/����ώ���:p� ��
 �\�v;^��p[M�!(o�Ha����Q�o%�ڣݪ0u�����:�c`p�� }cI'��%�[��H�fchZp�!Wi�$袇��d�L:���y}�o��v�HT��t�`�E�ǫ����3��&l=��B��d��jy"��U�n�.���1b?�����g��8�F* ���s�q�AZ2�ᱝy��z�գ�^r:-�`��_f\ݐ�������q�{RY𖣶LPM�ә��� mɗ�6�`��A�r�u��)�M��'�����wO�y����������#��F9�����m��麥�8ZOX��������'��)��t�8�ʫ��Ⱦ�%N�ۚ�#���Ǒ�T�~fc*����C艪�D�	yv9A%3eta�B���$�*���f��_Mgk���ȇ���dX��?xn%���n��}}�JĮ@���˱���{j����m`��� ��o)���E�0��z�-��T���~�,_`�^��W������iW�Qg2=T6)VSp������
lg6㤿�jj�̖+�^��Vs��'�$&J��72�y���\�D�<t/KT���+����jB;Ck�G�Αl
�_fcu���v�9��&-��϶	e��$5✖��$L\���i����D��[
�"HH�m�.��Nܶ^vS��Vh�IF�?���%nƌ3�,r���]�b���$�Lv�/�z���%��}v�m64/��`CT���]�g��A2�
�4=n&�"6:����G@N�3P�OK8z�]�U/�B�L�t���{%�0���VU��S��[a!�7�'�\�*�p��?�tJ�a`�ʦ�Ui�
���_^Rn��D���@�
o���y�x9�Z�X�MB�K���s�����	[�9�H�̹��_II����2�2\IO�����8�Ed�H�����E:Q8� ��+Og�P����JՅ�dP,��2ưR�a�$%wy0��ɖ��N�fq\j�e��ج�V(�*�����;��ӈԨf}����b�_/��}���&��&[KV����\�Nw:�:�-��d��@���( �$�3 $�m�Ǭ���ce36�/����ाy��m��Ն����5�[O����-*�uAͥ��')��xq��|��1�]���c��x�͡�Sz���dͅ�k�i� ���B˘*�^�%٘�����Xj�%uf��eY�ނ�J�$(3*uS�΄vM�߲ ��=�L����F���[�kwo�<g�]+�� ��,Me�XΠ�,�� ������re����[�K"댡�S��X@2�V=��r/M(Ć	��~.��So[C�l�y��C�]�����jR�KG�'�P�N��?���ȅ�Y��eOz*��-,M%"��`yx��rq�Ă"�I���~溭�t1bL�4�N��)D�+3Bz�u(����#���әԁ�����P�D�2�r&Fhoˌ�\�k[�o�:��,5d���ܗ����%1zo�I���I�D�	2"����� �����d �ujΟ��9Jl"puNYV.��8��8{�/�QT�j|6�`S�@*��e4���a����w��� -O�ix�)}���J�"JR^��݆����&|ŕ8�����a�NP����w}�ZL�^3ʗh�nĒ5$�3��l��D��Z���;~y)��t�B����CQ�iV͟�����-k#�8�AK�jo&��.D���!��-,���:���7���#Һ�C�}����Ż��U @�C|�¨O�g��Y���(�h���.���Ԗ6a��h~Vs49  b9�`B���J�7��'"�{�6�H%�zY6��u�I�yUL���|���Ȳ�U��c�pM9�7/���t��㧒���8C�3��`#x���߲�<��n�S[ 4 EY�N��S��h� ��M��;4Ň���>ix�����k�i���c�ݫ�ڛ�wh!�U�Sغ�u�!�o}���2�QXP�jǻ��1�����$f��|H��z�N��l�%�I�x�s�4��n,W�� E�a��/��ʟ�� �d��{�ad(]�!�m���`x�ks:n�޻�;g�P����lV}K7��s�CQ2��3��;�'^��"����foBG���r��0�j;fE����1@ �&�0I��Q����r��#�8w��vh���Vs h����=�2��%y�֚���׹ Щwų'�?y��JS� ��h��]��:��^�