XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������e\�}۩��;z��=��-J�K�y@x�X��+:(B��C��6^dQ���e^`���L�%@\�{�煙4�ťݽ���MI����f����{w'�lM�)��eD��S��z�[h��B%\"�m�q=$p���g�:���~U}��pd���`����3�:�hG�41JN�.�Ӛ	dy4Cqfׁ+-������{�NA]c�%�7�JS��O9!}"��*#w�_~�[��U��� ��c�D7�<�Aڶ��~��K�s��ë{qsk�*�8_@�닸wZ:��e�åf�W��y��P#Nxm[n23y6E���.�^\T�Q���Rդ؇K����8�$�Ί�i�T��Wm)��QQ�'Ul�<�p��l*U������ҀR��zk�"2U��<{`���3�j�s������L��_��hߒV���'�N<� &�>.�M0`�[�]�ɿ"Wj.���ַy5�R��-��Q�#�s�Bl �����}�<���4ʑ�NJ��Ҩɓ	m!�A���������˂������g#|�=v�ΈcW�j����2)\D�m ))ݘ�ؽ�ʁ<�q0%��w��1K�
�d	(g{cLЉ���Ȅ��U����)J=��b£T��r�C��`dR���豱�Dkd9�� �i
�Q2��>Ǝ����e�@�ə��P��*.�����7	ݸ��V/�pSY��8\3b�J����ۨ�Q��Ozf��;��]�a�@��j0�}o��)��rĴ��
XlxVHYEB    7738     790
�޻�z������jS�M&��(��LޞC��[
��B>��g�[��"��'�mm�`�Œ1�d��<5"�X����>��5�l1�@� ���D�������e��i|F�׷�N�x�K�6��R?�4O"���/8�<�8jaF5H�)�A�ai����"ψ]䀆�G� ���3�����ֺwg�������g�X�	��[-���}%�M��FD��c͢���I/��&��Ѡ�$=zi5/l��yG�Zd�G|��
��=l����x��<�۩)%�=�%�7ĵ��P}�g�
b!<�.��&�{�>#"C ���ld�F��6:����o!x=J�����t��5�����E���i�9�_��ʱ́�bj<&�a�����58BB����P����pcӼ��只�NOS��A�W`�����a��=��4�a>�8g��]bjН;��3-G��q��^f6-`Z2/��~yb����	��<Y�ƹ���4�%]�^�Q�)fME	o|pЏ:ڛ��i���aypv?s�B������K �i$��ɮ���@�J,�������wNY�A�3[��K����}�[�U}���AE%�`g���|-�mx�*E��49�;i�뿭ʿ،��aB�*�81O�:
�"П�q\�+&��k(��GۥN�n���!D\��E�^@���۱��,	nl��T��i_���RÌ�Y����C�Y�U�;3I�4�D��VT��):<tӖ������nLCW��T��24"Mtu"�@�tzY")�^�� ���i'�{=j8�)�}�>���lE��s����i�N��[���>�`���H��l�^�4�_5�Y��vǫ�~�'�V?��ߺ�4�X���=��c�?���p��.��
�>��M�����ѯ>�y}��d#iA�ϻ|�!�E�kb�m�&�-�-��V9$�3ƾ�i����D�J���rUr�m������%W�mr��e�aY �856N=\������n����f�I������R-KÚ��
|�*F�Y��Rz���x|J��S�2��)&�#u/�y���N.�K��O��%�Fu��^�[��РS�)��3ѩ�/�$�R������{���)�}"I�-p�%�8���l�к���� |9)���08�t�5-�����6�w�k�7�uI�,��z�mdtG�r����Q�^�����-����n������z�����b-4A�J	�_�dOh�4X����U��N�7��e��f��)#���Jm��;�y�,^���Cb$��~�k;�Q�,ۅ9G��UO��d����`���'j��&�Wb�k����x�>k5^�J>J��+�$�~:�t�����P�z��D{���x�]��d0��'2_AC̸]��n�I^l��Z�}8p����.K�GO�0�cN�s�g���|�{�����ʷd��L-��"X��'ea��NY���B�����m���8Y0WYZm��f�����	7�)�[q����>�\gl��@j���L.}�Ԧf8�fm�ԒLT�f�/zi��`&�fH�\��/V��0��QK�ύX���FA/�&3�����B(�/3#I���̎��*���qN�
��u�Y�'x���t�LBp-+K��_oS�_7ߨ"F�r�#X�6��J��W:I�f�C\��W�2y���98�bi?zq�-�&��O/��.Twح���B}��(,�+̣o�\�Y=0*5-���u7�ԧ>o�_�U��<#���͖Eب���ʠW�>a8%��2͖8
ގ0P�t�i�����I)r]T졦$(e"[p�Vџ�(�@��*!;��}�7�
W�\�ƞC��+&S��dA���B�D�*cQ�