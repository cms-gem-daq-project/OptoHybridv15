XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?@z�Q�5�����	�5�
�kc� Gt�ͱ8�B&#�N�~�Yyk���$�x�bҭ;���A����$6�7G?��i�k��h؁�K���$�PE��x����I�~�#B|�Q�F{��I��2�up���&��k��%r7���X�4��:y�wy?n�1O ��J#��������g�z|�S��}���%�+�n
���xbT�ʊ��7Iɪ�=�7����3!L�1�X��,���r}i���L%+�9����Ν���zA'PZ��}p�ͷ��1.�np��_����C	�o��O\�Eűp,͖�����\D��S)�$�9����}��3����M�5�?��
�x�m�J��f��iX�ģ(t��t}��U�rѱ^�'�X�I�{䣘�zM;����W7�To�ړѺ�e��r���F���i��-8�y�����?�M9�~�ϔ[[D{F�MD'=�"�!��D7��ZS����W	,oN�}w �Ҋ��x?)�r�)7�E���{����gĊUW�	�xp����BГgl���x��zQ�e���i�9e��k! �Hho�aF��g���p�)�S���g�HN�N�!1���`�����/��gh�%?[�C�3�X?��co��T9�6���V�|���df�8����+�!�m���'Me����M��%V�.::O�ԩ�F��07��U-�|D��K;D�3���xX���!����jkQ��ļ](�}	�#�HLP�
rXlxVHYEB    6fd8     c3024�?ґ�{v�2�p�#j����{�$Q��{����AJ�R��e��A;H��R��R����c�6�*�u|٥H��цU�'��3��9H�����s�:��6ڷ���=�P�[,��m\�B�H�$[�(0�&�R|���� �R�����\m
�qʴ�����_�(9B����K0��R�Uq1gz�� T������Gcf�%�\"~V�­42�1��z�ݣ����%�[K�S�MB��Er��_���H:��X=�|yHR��CM��=��y�}~�\dy��r��%�Rq�T�T�>���"r��J-�Ax ���W4l����"���ݜ��6�UWL@�׋{� +��+��J�.�."�[�nB@�W{���(�@yi:�ړY����;�k���� {S$�R���rS$n�ܪ�;a��~xઽ�X��~��޵����뒧��B��oLe���p�`�������K�/1�õk�T�*gw���q$$�828����b��}�W�7* ��s̎烛�p��`�'��q�۰�`o*狇��-��~	ԝ0O��ߑ�z���P��Z�hӒ��W阮e�W�|:C��z֛/x�{���{�t�9i̟W���`�Hg�pS�n}�śUo�7���Zo����S��|��X/��̢׈�W����Rk���r��ƶ܄����BK<.��{�Ԋ��x
k�>9�)V��;����u��!8������J�`�M��x�F�
0M ����!��V�ް"RA�M� �6�7`Ho;	`F����26��F!J�y��5���l�EjK�6�pTJk#ZR�bF�!�W�	M�ɂ��R'5�pf䲚1�)�ʗlre82)U�.C����m�e-�~�wu�Y��ӷU�j�h�'�"KC(�|��ԥ�=Q�HG�2s���Q"+��["���i��+g�d@�a�F|��a}����*z����Ã߇ŀC"�-9��(~#�٢_�<q�݉�/��27z����a\��)��_Q�ŕ�w�n �h� �r�I�0��oKY��֕��cW���e
�p�j��iǅ�B����W8��:c�A֏�t��q��WO�"n��)�ԋP+�]g4� ���A#j��@p2���ؑJ`ց_�7|<�Y��l��?�Be'C��f�﫩���u�o� /�ul�/� }�.γ�6���IB�c�4|�t�t��̮;�<�)�"����.��t�"V�bx�@�V*bN���aX�|�vO�6}��ރ�Z�u;h�dU�r|�l���O]��=!���7n/|��L�lMH��H��#���UG���1�ͯy��)����c���}i8�1���vm�N�z�z�3�F�8�#
���#u�Y��� ���C��������g��b��
O��F��7��sw`h,���$;���64��?���_��%��HB/9��?92��c4�P������"��a[�,�
�U�z��)o?òzh���ظm���@E��9��)dUb¬�}��	��Xu1�R���s���2�El�%�����+�\B�E�ݻ�30�ska����$z�Y|/�@Y �Z�z����Ǥ�+��(���q3��;��"���%�ʴ}��0Hb�>����p�dh�~��t��Z�Z1�r[��;���Q+��F��[���J���Ȳ}MD*�/I�!w�b�l��s�����ݧ �U΂���B@�OX��ޙ�����%x]�7�ʛ�Ld%1Y�Bs�=����S���Yqq�@i�V΢|���Y��5͹ȄXB�Y�2�|=5!�S����6GJ�����N���ӵ�Z\�zPm�f�����%����.���b�7��5�Yi(a)V�5S��BG�f�(��Lر`��i��1m���<�ǏA�2;�m��u@3��v.'J�p�.=I��ļci���z8���%m��>Y�:�z�aŷiO�p��������wv����"au"� �;D�L� ��}~�õ֏��<#���6�e?��2L�~W�����ƞ!\��n]�>@}�r��z�!��N&���pq���Fs�j�7�����7��D�l�}Yp����N�7�ij�/FD��P��,S.nyXvXjߝ�+-d�K��	�y�n�߿	QW�7D^�D�9�߿;J �g5'��/�Mԫ	���R0w:Ons��*��!��o�z�����kE5B��o�Ba�eB���Sbo�rB�]��wz���?j%�SwK������c����O�k�=�kl��'�b�S�	�g���bG��G-����O1o*�&�jiJ/� �X,��D!���7���:��0��D�C��<S����6f�h�r'�� �3h6̓WR� C��l�B�/��ݖ�	�˦��)-�1V$>�(lϥ���S:c�t_��]�O���Jv"���!� v@�½_��9���v���">��*pO���B^b�P�8z������Q{{�zY0���!Y7���K��m� �u�
��2_#�Ԛ���I�o��;&`1��B
��g.��~����s�!6":<Seヾ+����������W/����8�A,>�q\��'�rz \���*z��h�O�f��M*O��3[�E�E��F��$e�|L�x�� 5J���^Ӹr[ᰠ���Ωu:?�9%�U��ȥ�+�J�%Tdl��-o��*J6�����L��\D�z�z�BmBm�N0��.� �a�J����&����k��Ċ�o�0M �\�"$b�n����K�ī�)�����mi��N�{��W'79��v�ω��F���c��ۑ��,��4��y݄����5 ��mi{'�����vK�;�a�q��癔�d��z�d��o-��4d��ǚ�ThX�.e�֋Ʃ�G.S�2����>97?�o�i��r��y7v�ؚ!�<d�3%5��ȍ�5�D�V;o#X�;��62CG���iwgQŊ1R��L�����2G��=n�n_�V9�R�0�^BI���>s�����=ah=�Efn'*�92��W�+���/7��dq�i�P�bѬ��qn7���*�I�:2A��ͳ_"&E���w#�D