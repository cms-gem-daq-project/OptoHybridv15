XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t�(��PD��6Z �1}���/#?බ��̢B�����sIϓv�йe	5�}H�K���3C��q�-������=�`}I�J�.�3L�gh�,��]~7��hj���#���쪒[��O���λ'Z�{�ę1�k���c��<�8�M"0xT*��Sq�45����v�+�j�65&EjJ+e�WN������ B������s��O�R�3<"z�H�D�2;;AO ��@����Q+��K��Ubގ�f�_�&����[���Ɲ�0�P8�|�|����=11�;u�H��0�y�&?'�SQ��K�m7q�y��Ԅ6�ٺ�S�jGP��F�F�f~���c+��$�r�^��dAl��R����@�cՀƕo�&�M�F�g��MJ�#�'�Y�4�.����k&q�K���/�Y�WM2��5���'?���=�m�a#gݶB�?.�����;
}�����{�$�D�^BEs�)�s*�<˽k��V��6��v���q�>�VZ��r䐈�=�8�s:G��?(����?Z�_��N�l��c��p���=�K��qT�kg�c��j�p�cE&w�n}w���%g���Ж�y�zz0�qL9+�_�f�x�=����ƭ�����0����d���/ţW���l�7E���2�����=�R:9��^4���,u/>3��<�}hN=r�_8I�Y��
s�:x����g ��BRa��(�b�����`��I�!��Yt:��l�^XlxVHYEB    50aa     790����vM�i��Q���cR�����������_�xLQ6z���|�>L�D��笹�pE}��^uf�ͷ9"���z��NĨ�x��M��olL�����S�{��/c����V:��hj�/;(/\(���*�B*���}��(Fߧ�}� �ѩxY�[��A4Be�벂��>�G�<R�H`ѫ{���8�W�eF&v7��5��Q�9o x�˱y%Vk�F2A��ѓ�#�4�X�=n���t��;!p'ѵ�i�X�?����������dNNpN�U}���{\��:�?N��J�D�D�'�T��<`�O�ed�?%���\K��㩳���e#���*(q��V#:�Oޢ��X@L�-y?Z�9o�|Hv{޵Q�M��;���L@�LZ����ӛ�(k���T���&mfv�]�/$:���NK>������F�O�$%��	�o� ��zLM
��ݖ9�� ��	�0�����p#�!P��U�'�-�]c�ӈ��S�z����qɅ�1�P�
���=ov�_�Xܤ7��%w�J�qK�(�l��\�̑a����U�v/�Oܺ��q�՗��g9��&�������0�-l���!$6�fhQ%_�3����v��|��017ğ}q�˹��Ig�}�eC��������=B�$���vS[Q���U9\�)�+y#�%�p�}D9>9Y�Hy�DL����'2v��P�0#�sj�g��"��k_��91�̑���?�U�V\�L�[��[9�U���*:���Ƹ�#�7M7;��Dbe4�,\�؏���߄�y�sþ��7"�J��wb��}}�O�^�����z&:*%�cG�$����3dv':9GJ���|�
���]6��]�1����c�DDw���p�%�d�X�׌�'��k3�i��{o��,���:y������Pڣ�K��KL�ެg�cb���ǵ�R�:��p��¦��ZИ\B�D�����Ȣ;q�d�������*��kz�ڞ|TX�nm3I|�����d�^��������eޞ�0�I���ڄA��=��� ����k�#_�ka����ArD�A@�U��j'�q�M�㯛�`j:R?��?�Y�F-�ً��j
q�U �j�j��,�#��%��%L�8�?
�/�Śp��O%V:Z�
��c�\�� 2�����MN	#y�V�Z�uǸ���0o�k��ƿ���lg�Ta)�W�̔����;|P?R�˴���Tމ������u9ʰ�:�g4g��I��r_�6E�sB��w�Z*�#�p���� ��>.�E8}v5ќ�7������L׭��r5��(��kl����Z:#x}7ۖ��2������vsB��~J]���s��o0a�P׾qw�5��!��w^f$+�T�	Q��HLx�ɦ7�f\�.e��?��k.}(� �>��$�f��#������(��K�Ϫ�.��Ւ(]�ݲ���t���8�@pR�,�Z���B���g�8�����2�B�[�}H@}�a È��{��R?��Gׯ�s�a��OD�A�g�Z��3���Z�+�''�&:�������xj���R���藗��#�ყy)�8�l5�9Z|��@�[�n{��K�W�vz����Ӯߋ|r��4��+8�X��/q8�Kܐ���������ê�{δ�i��"㗫F{@""���~.B�>U�i�
;�,.����k���kڣ���X�a�,���t�i�����[N�Z�Y�8��^%t ����՟p�����1W�_}��z�n�R�R��+�l���7<T���X��I��=[?�E�B��RõfW�dm��e��M:c-]H��jTIb�w���/��L̒��qs
�~ 
+hH?;�F�����C'l*��[��eu�'��:�!�Em%�