XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U5��/56��C�g�����"�����+���qq-�L�z|����=*�i,J����%V�hƹ�T���b�k��& %*-ې�L���[�z��x�Bs��2Y?�prR�P���|GX �N|��=K���Mvd����I-"VU���+֢=���s5e�gn�*��W����U�E���!3������iz�X{��7V���]���+��	�u��Ɨ+j�~-���N TU�k�u���<��Ul�8ސڶ��d��! ��H?}��p͛�\pXq)��!`H	OV����Qq��%�>��6��:�ه7�>h�Q9�z�z�*l1�A�X�u��H������=�����hw��}IB�~햰�J�Q�vL�����n�;l�M���� 1�����x���o��Js^����������v�G��7Q��]uq>�k~0�#{�=�@0<B����M���?�V�)=����L��4�������SV(���Tܮ�GQ�0�'����]��� �	�8�5�b-��Ŀ�pU9� �yR���n ]�J����A����34�0�z�|IV[��$��8f9�E��%7�&XkL��� @�����G]�2��ܮ�%� R���?�}L0���n���bh�Ǌ���RI���>ʄ�ٹn�vrFX�<=�=X�e�\�:��yj�QyP��,���á���l�i�����fv�4� 3�T���&�����0բ���$t�ʁ���CJMm+�(4�)�m� XlxVHYEB    3a1b     d40�r3�i��&G(�.Nk����������' �>?rq޿���X�RX���e���_Ea��V�������M���s�o�0�G4<�8��j ^�"�i'D.��s���L8u��y�eMy��gicY+2�>�p�3+�I3��Z��/��|��[*���(vŎ�}|8wH�M�ۏz�0�y�yq���(���d?iK�Qj��VI�U ��/b<QK9�eL4
�����7s�G�X��q�$�D�5R�������0��a��S��uM����T����6\�R��,�poj�¿-P����(NM��ώ�E����vmnO'��>�9@�2X^b��xY�t`
m�@ ��f��}b��!3�ƄЗc�,T��Sk�i@����Ʌ��P���T�<i��!>B4��-=�G�nC�����V:bX�Li�`y�)�� 7ٖ��ў��S����Mj_�ؕ�r F���*�t�-��ked�dnjB��?o) Z�<��q�=�͎d��`�K�"��Eo��rQ��������*Is�p"se��.6!Ȏs�>6�=d��6u�I�S�%�eJ�!汎 ��m�� ��\
�6-�<���:�߳<�T��Ka�{�m�d�9��N� /���?�
���]Y������?U7Hb�
�E��XI1��q�>�M��A\����L��<�:�CL��T��n���r���D?3k��� B��El+Ĭj�ʯ��?O�+��g���5�,1�3�o9*��7�$��I��P�u�Q:`d�¿Wu��>�U�55�&�?*6z��˸%��!��<R_zP�n��45&��")�E�
���9���y��\a�B!Z���N(���5<�WXW�����0R2y1�ڻ�]�#�A�-3P��FV.�Ӳ&������c��E�'e�KC�)1;��0/�v�%\371ܩ�=��Z7�4� 
��:J^<����j�<0�_���u	ka̝7'���2
j�V�wj�����XRM����d'�Q�)�^�*g:;����k�)G�h dp��O�M�����v˗B w��6͹���������y�g�쐇n��M��Z�[yl�	oH\�b�1��za
ñP`/��1ŷ����
��T(�dϗ��C��p�d�d���Qf�~�ek@���Cu��[�.6q.	�ˈ�������]A�"�zc��`I(���	���ǣCK���Q<�[1���S��wP��������AU,�C8(�D��Ɂ	ñ�qa��"�A�lv���	ϔ��$x烶A�>��z�;:`:��r}��k�H�A�ym�r���oB���ߢ��eo�]r0�mf�nA�l7�%�/e$���VڎK63�j�+���s��T���������l��K5�'��5[D�Ū4�Q����K+��10�~և9N���C���ܻ�Y�6X�,��H�dK~k�?�)��aG�5����W+±2j0n*rS�h&�ë�Vm3���}�(�,��a��t�ոW>ʇ.u�	���}��"9埼���tC�3g�@�s6mO�%���T�.l��v�0 �F��O�0���)�B~AL7[�+߷�t�C�͑���pA�R�"L;�D[葓�ݥ�q*'��g�.��b?:��a�Η�znvgE]���=�WCP�9��La�1s����i��#8|�q�h�_���b`���Q@3��I��]!�
��M��U˙�,"��!gO'N��2�4�B��2d~=)�Q��09` :(�����^*\�s�yف*���4l^�ᅂB�ii����x�`�j�\@�eM�>�ע^�㽇k�΂�����N 0#Ѿ��B��%�~2C3���&��[��ќ#X�l�}]����کXh��������4(���2��l௦�ebC�@c!p�#yn+bVJ��5��4w��Pϧ��$���G�D*��֗E��I� ���V38��*r�7`�P������v}^؈�qqy��ϨYY��C�d��u���l�_O׼��S�H�=�<At��s�J=�Z�Rx3�Zh`�~���xH�}�3K�#;It��b�֏[���$���P��
EY[5,t>��e/U�����}RT��磟����=�ۤSOe�
�$H->�z��r����4&���7�����%B�G\m�����TP�Ž��FJ:���^H���XY�T�<͆4̸����ge7������qsp(<�E24���yy����ޖ��$@�����F��b�I*-!J������^����ܹ	d��C�l�Z̈dז�U0�r��}͜Z�G���%��+H�@*"u�~)SN���In�>k7d��!wM��+�Z�.r���]i�ʏ$���H?e���h=�؎��[ҕzX|)�=��]=Z�;�t��)����0�d5D���
����ZX��e� �@�D�o�S�2�l{7,e�[H���˛̑dР{LmN;>�hb����Y��ٻ�y�};��G��_���Q���	8-�y����2dU�4XB�6N$��x��r*V��2���A�PV�W� �]��K�l�_�-E�JSL�[�yw�9sL�l��[�4��,�,eA��ч};f�ι���%~��Z�:l4}4N~~	�l3��6 E�H�k����֫G:5��в�1�_,��L�R r��~/��8`4~��X	��M���[�C;�~*A�q����:�@��^�7se
4�Z�:�9�kR��١��Θ��,t4՛wC$6hōгV�1RJsk���V;s�w3���sZ�D�X���&t��w�^Z�/��3wP��y��{Ǖ�n�2��'�[Zƛ�ay{~�8l �Ln�說�:��b����7s��}��K���e�֧��M���0��
2 ��t������wo�n
�bJ˥���1��s��2W(i��	
9�fz6�C�z�e2����$�?V��c����z��MK=a��)�E�OMP��_F���ٴwb��J\���s�͕5B�+��G6���>a�l��w@9��,���HY�F;-0�z���o�a�Y�O�$��U�:3��m�+B��u/v�T9 b�]��p�i��t6������]�q�T@�?�[д�.��_)��N`�G��/�e.nI;U��Ч��S䱾[����MR�Ӵ[������;p��x b���RM��:7��YzX$I�PY��Z6�H;(S#J�v�|��b �����z��M ����D�����oO�{\��PC���f�˪e4d-~�D~�R4���'�oH3>��f���T�	��QX�cø�u�p9��/�