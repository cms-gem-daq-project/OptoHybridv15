XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t2�|�?,�:0�V�]�der�`����U>�'ޣ?�z�D��/��w��˅C?�e@�)�Jg�ŀ굮'y_�D�È.w" �=��yKӏ�>��{h�>Uџ?j,�$e��j�.ii�f3�����(���:;^Ƀb������������4���4�S� $��XɖAE
A	�0�=BVW��\�Y��B^������}
�/w�ݜC[��d����W�,G�w]YF">@��g3j+B�����"�m���ob�%NT%�=���9��{דlӞ�A��A4xrd8rZ���	v��ZE���k&�x2�zR�_XȘx1^T��If�%�i~�:�v6�_�Z�K����T2�P��t �1�_�D"ͤH�@3e��qS�o�c��H�\V��;�?����U6N��͜���.�@�і��=}�Y\�cmu�����b�9
ޟ�cR �p�W$�ϸ�X#��λ��.�N�]㇈a�
D�_"ڎT��M�r��9U�˂!���/��Z��cV�{��>��\��ǰ9��B(��y�\�[�u`Hn���HhF{	��%#�*Ә�u�eMF<c�l���zI{1�N�nj9�}յp��o�O��%p�����Br�w������d�x� ��AN~y;�1|~�Q�]�>7p4��J�^ο�<r�vI"]������#��^�ݼ�4v�p&O��i��mZ����:7���	(*����#COsP��ۦh+=��m��&��{XlxVHYEB     bbb     480"<�A\m?&B���M��3�k@oG��; �K��M�$"�֪}N �� ;�?�	%r���_�y��-B�z92U�M����8���A72-�ԘV}��[H��JD����� P�{'^0�'�@H�oR�e�my�k�N�Mx��qɳ��c��gu����'���8w�|`k3Qd�~D��������܆�k�r���V�!l�X))$:�~�	��R��&��@�&�u���Mx�:>������$���w�^p�`�6��r����;E���7�aA	q���[��͒1͜O~I�;���5@� Xʐb����Se��������4�h�����p�P�rnU:�t�3���E��JɁ����'�:#� BFh1��y�KoΨ���H}��F���@��N`_��#�=��6�gEw�'�	(�,QYx���Uh�\�6;䁨��Of���y��7����55Y�j��?C:��, ^}L� '��#7l'C���븞����-g4r��_�<N��c����<�N�"���� �<wC�)���;�U�a�t`z��%M&��O�s��*8&[�P��J�_Du���cX���*����^�RY��)��"��
�Ͷy��r�~����-�)OD����3�OL��?��n� 檐�u/�����|�M�hu��_d�%�O4�H��N�J��<C���S"{��`'N�<�Y����� Q��\ϣcXq�sI���~��Ck���3��L��,,n+	������Ké���f�ی�_9�3�z���32]�FnL��%�-�'W;���J:uY%�(�yw�n.�T(�=o��x.ɦ�X�L��%��˗42�.��[(�ׁ:t_gx�O�YJ�J]���4�~�O+��<�aP�����S��|uށ��{�Z�r��8sP2�{i��j��PԿ�����9�{��H	lv�J6��LN�XK��r "-o�E6��[���k&2�[�/��L�f�O/G~̕�tNQ�qzM�>ЋL�Z��n+jd�[�>�;L��xD4�C�l������[�@tC�x�͏YL��
��Aj�^�W��20�8��U��+�	& �hG�<�W���D,�Z����b�������������<�?