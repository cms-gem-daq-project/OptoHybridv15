XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����9��Y�����8�~!�;������"�؄E;y˖�X�=A�4Rui�]$�u�kШ�".߀�azl�E��{�-�#��LT�jz��ct"'1�.�Z�[�
gW@�HVݷ���;���������&����h}�US
H<3���e�-%��1��x�ܢ�Xbh��3�I�(���~����
`m1��@���y3�ŔT�M'	(^[=}���yiM'J�	)�79N�v��^��������5$�~��m���A^�Lz&�F�)e�Ff)Z�㖋�DNFHU�,t��G�!��Iӑ�� 'D���:y�jvTҰ16�yp�L��^_q��:z�>��j�H�F#rvf���2U��ҍ� �� L�޵��ݾĀZM�g�@-���9T�1?���ny�����@!FK.���C1�ܳp�[����Ғs�4O��P��di%d�#�7-���i�q������Ӳ��R��W�-�h#ZX��\HEbT54+�R�("�pӚг���z����H!�����;�Z�a&�v?�s/��m�XK\Α��2¡t��U���j���O�7�R�4��
N5�`����"<;K�E��U-BB'��M�0@�P�!J�3:�?	j���!�����%h��өE���"�n�ʉ��+p(2�S���)��\mu�a��}�+9�j�a�UAL&�Å�e�F��L����1�"��Wf�)
=fkՑ�A�n9jՔ�Z(kb����� QQP�O^
�]�|�	w^XlxVHYEB     a3a     370�$Il\���k/���5 AZbŪ�鴤��5�c��Eb���!�|��@D<�J���p��E^�X=�
�. �f���푎��n��$��+���e��ݾ��R%��v�7����b_�ĝ��:�% \�tHb��pV���v}�g��
�l���_���Ԛ�[���n`��6�l�<���YG*�SS�΋rP���7����/�F����^��e`�� q����{V����������и�����z����a$�Ҟ ,J�
wBA��|�~�����~��uq������!��M\Dd���F��̖��t3@�^[�L�LT�t�vw|�E��H� SC���$TP��D�s<����L�!+��>�6���m����0�˗��i��!eǼ (a|����9����Sٮ��F��7d��֜�F�Z�<���i�F�����|�tҖ��i���ԏ,�j�����t�j
T\�:�bꨦ����6�y�;T�- |0��qz��Ԥ���������V��v3;��mX.W�/��t�ߦ����	�VVd��ը������g�ђK̍P�����_l�� ����Z�R���xa~UT�v�F�����b69+������ͪŵ���;�-x21��n&���Z\3=�ү�<`�s?��\�m�!-�Y�b8)'E�p5�ҞaD�3��7�x�0�e� ���|*�2�_�u�; t6`�y�wF"�^`x���h����꺗�Rv���rLf�]������}*|j�;��J|����n��*D�	M��dbyj��L���%ٰ�rBؐ�	�1��j|2���<n�2nᒶ��z��@�z�$E�