XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�7Ң��D��H&[���������e� l3rFB�P_���e�9z$?�6EfH���[���U|cT�;�:�,���Z�+D帵�/������Z��ʓ*g���B���_�9S�|��Ռ�gfV�-�%F���c�r�r��>���~LޢJNH��!�;��4�t���~[�2����d_��+:��&`������l-Q���2�P�M[�e� F��B#q�W~O��qKrk�����`
jQ������+�6�4��Jo���">�$o7'�&/���Jzj�����@���MT�/�°�̜�=���X�
ٶwq�9�F�#��q]\$��P5�C?�I�w�/{A��yJ�.w��5�|A%߫}�,2�7Ԫ�*PL�2<,�`���~=+K��DH~f"�86�Ye�����"D�9�5)~%ŗj�����,_p)���A��Qx���f1��&y�w!�a^���O�V
� s��e�b����e��Dz����{���N	��k�p��l��xQ������f.x��[�M�S��Hz*z�<��_�rs��5��q�}�\�_=���u:��Z(L3� ���^ě],f	�Ǌ##�R��N6�ƌ	�M��2��;����uF��=|SD�*����B�/ު�.��]� ��ʕRpu� ��9+B��'�Fˑ���J��m���đT}�z��*�ګ��$"�=��[b�Zp�,OO�-D��G���B�Q�-�X���_�&�ɛ`s���m��/�XlxVHYEB    4d93     cb0#b��_��k�h�ZH�,-�.��H�4�i19��P� -�I�E%`��aM��A��<n�]��牋�	��SN�!@9�jǰS?�x9����E���,6R��:P�b0��L*�Y��C�y��4�a1���qW��q�B�W���r���J8K��y[�'�����*5"��#�a�t��d˸��c��y�цb�#kp�}��v�/Eh��*G�FzJ*X�M����b�=�w�q�89�.����\���>�r4��&�ˌ2<�8-��֥��%e��L@0SK�i�]�K�Wv�Ew�|���"��p��=��αl䞃&kw\B*�x���I2��7�z��]�*
:����}��{I�x\%~�;��p���@B�s�N���<��P~B_���\���7�p��	�"��61��yJ{`�v�"ú�t�	P��$ Vp<�����+�܉C�3IÂY#�?�B�#lHf���nA
�m7�K�F�R�`ǘY�I*��x�b��(U7�" 
�Wi�B1ޟ?�sYFF�K	�*�^�����V� `e�)N��YG�k��:dڻv�3�>.�ÏKm�Q3Бs�nAU>1A��g��[ N��]�� ��O�c�NJZ��� V��,�h��]F�W�mXD��G�f(~g���o$`D!Qa������$�p�R�rZ>��Ң�{���\���G�.�wfQ�8ju��b|xW��]U�_:b�J깼.����-]�[���m�A'�4��8>҈�[9"�p�M����'�����+�D� !�S�G�hv�p�P�fNr�3���ЖD�;��h�t��xb����}xSF��ʱ���_���$wR��!�����Nk5���O�]NB�_���\H�m��c�hȽ<?�i.���W\F~_��A
���Y7P֮Ra�ףAf&a�����T��f9���`�j���:.���[������*G��/�N�Ҩ��嬡X�xpEkc ꩅ�ݖ�É��U>��,������E�)uG�zkG{	�@tl��	OW�+�T.��H}OYxfU5ה�������ǆT7Nb�1���Wy{����0u��f��M
�{��x���z�o�X����fv���`t���LhZ�}����+��;,�γy���ڄ*���ij���L��>���{O�ܵ[�+	�qyWCd/�?��J�?)2\/��G��ȥu`�b����-�j ɨ���Oc�s�����B�M�M�_=W�Z� ���������*��}��Dj�d�R�����y�,�& v'v%ˎ�\9I�[#���j�����Ez�x7�1tW��9X�7�œ�ؾ_(s��׃\kqȣ)7��gZ�a�0�c�r������\)]�fs<�{0��h,�&��ێ�(rp���0��b%fᠻ����炕V3�3�/�'Q�ۢ���ڲ%�	��p���6�(GXf���Pg7O��0,DD��U�2��f^�vD�.>��!<��|6ĿpY��vHm�XŌ-���3&��"��tp0AZh��b״�&�W�8��]	�]Nu!J v����_��Af�i�Y֙e(TU1D:�-��>4�AnH]{�����z��W��]OLu�w���=���66G�O�yQ��������V*Cr?����s���ܾ��"�']���n3��`�jH��s��3�,�8����e6���}k�a$��nd�O)���oݛ��h����K��`N�+ϲr��4�;Nr�2�	�J����ŀ;�s��c��>!�Wu�v�)����5�6�3���hS���L��1�WNhR�]���� ��f��F�40���6U	}�v��+`!���r`^v�oP���NYy�t��մ͞�a���m��D7����5��n �V�x��������-��eNh_.q��%+�ؽ{��Ȟ�β`r�Ӻ�\��xáqC)�@ވ��nQ@�>�P��s�'����,�|4
4�V[��#�c�f�i;S�b�� q�G�5�z+p�vN�7�;ʫTU��~U��v{Ȟ�����Y�%�׉�� #�(�Q~!$�΢�`/��48�Q s���X�^��V'V�!�+�[d���%ͶZ���a��;��ݜ�\a��ʺ;�c��W�Sۙcِ�<q{E��y���#o[۳�W7?;�@$�V���>De񏞱�����?SE����A/��������E�j#ď��C�v�=F���r#&g��Y�u�J����V��E�}�8�����㉧өƛ1L�����i,�G����j����+{@1�����# Y*]6�E��vnux�ϺQ
h�rX#�ӫ�X�ҿ쥮`W�^ � V��[G�3���v����a�1ײ :�5i���Lh+�v6b9)e:/!�����d
NWT��-���U����%,����Yy���[@-EY�k�.�V�@�"fJi��XB�yֳ�Ey�2�N��l�������UT&�U}[��Ռ�_1t���39$�n$�Mn����^�9���$���f޳�Ub�!���9W���O�!���[�4��ĸJB��YW�=ۡ��P��D�=��S����^����%E��Ք⎥��79Ӈ�ˌ��*��5���� 9r:����r��.�F�-< !�^�ӚuSu:��O���?����UB�,�.��~��e�#:��^�h �6S��@n�����}�`NRv���;��2:�sX(N={	x��,��A�/9r!(�G��~8.<k(�]���>�&��^]�E���*�gz�Fc~����Z�߆�qHQ+�#���R���J���K�Ϛ�m��ĕ�xx�}�>�(b!�D���V"C�����{�g�/E�
�tup+�V:�#���]g�int��p���Tl�/'>�8V���aȺ�����"�r7�1jP$r���U뚝�5��������!y�cmI���"����6Z0�RE4�˛�����s�S?��El{h%I�E>���X/ vj7�}Z�`�4n�EUf�����s���*T8=P�~!�Q�@q���O�����ٌ�iz��
SZ��U6z��,�<x+����
�#9j�V�f���{���x \c��Lg �{<C����j��<�-���xt�)< �"eIq���+˺��}�(2w�Z�P�i�c