XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ge�����Wc����pG����T ;�tk�y��}�����/��u=dA�#].!T�Ih�pD��a{�?f͒q�&�R�r����Gk��Z���x���&׏ސ1����;&3��&��p������}8�5�;�:'��Z�F�1cj�'2��h�[];�о�E�q	H���c�?��57HH ii�d1l(^�6��A�`NZ��y Y�ǂ�:��{2\��A͖���זO��c��{�"��.�:���v�ߦ��[q��|*��B�A2ւ�7���u#��� wof2�H��u�l+y�)X{�yJ.����6)jg���E���F� ���x��ڬ�t�lUč��r�c��Ǝ�,��N�������#���X�}oKH���BNE������`����9��)����eu��9"����󗀿'��}������A�P��cg���=���	�y�U�1|��Wn�|H����Fߋ6Eѥ���BK����<�D�7BJs-2\�J�����BA"6�5iÏ_��]xO�"-��8U(�-�A�g,�sJ��2���h���O��i��`L�>c&e�J��7�����|����)�߇ij7�����Z����ϫLޱ&�a.����#-���������/G�~�(����^<��[QePL���&-u�9�����):���cm9!_x�	�8t��FR���S7u���7��\��r��6sXYъ��+��:;��!?XlxVHYEB    1f8a     780�M1c,8Jұ�o�����&��JHd#V��;y���R:�{��Bx�����������븦����CM�
zpϙoMwi�#c�MM6�㨔[����W�������D}}��� �r��+�U����cs��)���s�ކ�?�CCxZE�m#��($���9v(g"i� ��Xn��R��@�|sgީ��ƙE�@æa���v;Ȅ�c���r,f�|W�Y�[j�Pդ��'�J�	&¼j���D����JҸ�s�~�f4��n�� F�{�"���,��h,��N2(!�Ȇˁ�*x�%~��ň��Hgo�,U�I=T�R"Q�!`���ǃr��(�����̷��I����\�������H���H>�
pu�;|uo=��̟�jn9[O����x���Rc����>g�F�F��#�ˊs����W0��|vl�~�O3���ez�v �ok篞C}5�J���Უu���g9�����6�l�44���Hm�y'��C�%��c�b����kֶoi��
O���z��1iMP�V�۶��������Z|�}���x�$�f�*�u%��<%^%O���K�]pD�\⎛�=�(r���Xp<�
�a����Ky����T��M)������Ҷ����>���j֞e����AQ����t���m_`�6����{�W6�@AB ���@I�[M�[	��,+Y��_0������:��sD����z��^m��Vh����	�>*�ˁ��I��dq�� �[����%J�/�apQ_���H�ٌ�^��,5�A������AV�1����i}h$��CG����i8���	*�{ZϘۖhxZ�Eg5���AϬ8����"E�yJ-s��^�Z�Xm�T�uL�������;q�"}>�<O�Z��F����:��T��M�^��⬯�魛��䊀;��*�q�ϲo���g�t��ݷ g.�{���ѶJ,�������ˣWAk�>����9�8p=,-�eB�_���5q+h�|GB��53��,+J�¨[��.�oU��'�	U�3��&���/��2,ӣg�krॼN����l���C�+��b(B�*ړp����:�q�ؘԼota��Q�Cc&�%U�[Ft�t�H�KN�@���r?/E_�Q8�lH�Z����޹(�*�|<&��L��%�����V�aN}&k3"Sg2-��N$m���&�°�($7(*��Խ-⏦s��힏��=���#ޜ΄��l�� ���Ⱥjͽ�x�@<�(�S�� ���L�>^.4��D������1�ݒ	 ���'��p�G�$q�:X��c�@C�47T>]��K+aR2RqRk���ռ�!H��{���LP-�:�ƞ�Ά,|n=��X/ĵ-�ˎo�)bԲ�׋�eug�պ��^8�.[�=�`��b�2���J�{�xn��BM���v���i��?fweiv��n����m�f��~�_�=Uoe��>��֩��֩l�)h��$S�zv���K8VYB>��j �Gl�#�S෕����%��h7��^�L7O��:\fH;����r�/�a�~�%6x/7�ȣ{^�o�p��1��P���طe����Nۿ�W�аFU��Jʱ�M��U�4p�`P��!/=��T��M�TI�9&�Jo�����?���&ң��#�����`��K�� 1H؁
G\��\$�,Ϡ� M�!�i�!�]D�z)�0	_o؋c�</!�К��a�f��ᜉ��ސW%2^�U�I��e:�����P�J·�Nl53,ؤ�|:�6)�^�W�8Q����_�jC8���p�3�:��J5x	��5F�O�f��~PG�,uI�	�^)�ڂ�V�g��