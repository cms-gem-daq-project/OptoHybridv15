XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w���M�~	�?� Bs/�!�tP}xa�4��:Ch���������������6Z�p��w��X,�hU3 �G�G��U�F�r#��3�����|x[�C��X5�	#��k��/w�bA}���8���W�g��������䡳�5�(��vw���WE��ɞ!1A�{q#�mHȩjY���Y}�o����=E6�eq��BanK �Rd8��L�C�,A'����&��(� u��?K�H#�:�L
,������E�2�X��0����q��g�`m2�1@��d�3fĤ�Ru�K����n�i�����1hR��g��^&���'�T������X��{<|�,\��O�z�B�c ��D;�������#�_
WvC�Y��	���OjZ�Å��x�##�����*����M5�s�븾� ����3E�"����]0`�+��m�����e
�����Y�&��6��5to��}7!��8ðX��;�J,y�I��u~6�h��/��L�d
~�i��?���m���-S͘/�l����m���D �X$"� u� �~el��U���a�>9�01�B~Cn���9]3i|U��}�PE���%I�y�KH������)D���0D�RI��ik���w����ƥ �x�nTg.�/\�{) ��c�����B�<��j����钋z~HCTN|��pYp���,z���w}�Ck��c�8�%��0������'�x���M\l8OY��?����؄�)e?��XlxVHYEB    10b5     410lN��M9>�WF������*wmP��N��G�EӾ���[T����F���	�oo�s��pW<��Cu���o���龃N�
ь�e�P�.Hz"�T�'�x` �#����R�]�Ot1>��r�ƾr���X���3��[�=`��[�ۧ���J��K�f��G��,�)�D� ��M�� =�4K�>� � �� ����x�~>y���$��џ�����1��V�����'��Ad��mg�<�u}�b�d4�od���ʃ����(M�G/[���S����v77�'d=�_A}��c�k�\�JHh�/�����Pw���r7D+�i��7p�2G��u��h�zo�����^����;�vm�^/���<��¯�7ܯ��Q�݉~�;���i6�Y�M�Wȶ+�i4�8����$|��/�.Π4��(��߉d�3J"�]
� 4��ztJb:
��h��3v?+܃*\�>q�ߞ�4Y�ڛB�⡜sI��Y�A�j��y�*�D�Y�}��y`Z\U���аk֤�P������RJ����>�~2W�<��iَH��>'H�,�i�04��+��`e��]?�*�'zk���Uï�2N���h�Zs��
�~��?���`�*gr%�p����j��HH�uv:L%���pa�Ud+��Վ����&��
�j���������%�Jȵ��J�t2�y������p(��N���Ʈ���ڴ�l���7R��Y��=y�xPw�D8�=e�V^M�(���l����N�_E�8�!�Qw8�_�%�1]s� �G(�@M�o�*p ���s��}��
#�ߤ�G���(g�`�6��繺�"�`
�����^G�
̓U6��"i��=Ϲ<[0���z%o��9���-7��?2__��@c�]}��,B��4"�D�vrrX����r�֠y,^����,_Α�:����q�}71t��,�ߧJp��RP����f|�
�L�]2G� ڧ� �2��d��v�x��o�0�?����5GUk#