XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4���?m#��JW�8�\RRPk�=���I��.߽C�w�n��=�(�-Bv��* �o�!�,�"���wK_|�Nu�h:^^2���~���+�І�V���	sc*H�]*�8҈��m�C�OĒ}��u� $5�6-Ӿ�� ��b���9��աeǺ���L�}� x�,���ǑT�դ�OЀ�ŷ�b���}�v���Wn�Gj��v����z\�92�����o<Q5b����g�S��0�}Hv�w�LU)�:�TXo�H���t��P�NX����(E*���fv��f�7sJxv$Ѷ�;�'%�(28j$�������c�j(6�����V���[��,�1��d}��f�肁�_��`��3+&@'��!�CҤ�ZЛw�-�㽽�\�@���k�G@�X�������ۿ��>�Jŵ���^{@���.��7��d4�ȅ���Z�`p�%ܑZ�y1�f(�P��S/�w8�D���j9>֗�)my��HCs�O�/z��S�O�]mkj�y3�TYy�ӑ����Ag�H�5�q3TWk�
�5�2�+	�م��@QklK�q �'?�P$#��o�",�Tb��;0����@t�m�:��]�WGgA'jZ�/6���AU��m���E�.�/��m�)�yO�^�ƩL+H]@dG��^�;�\`�F�V�@���:F���-O��9�|��i�:r�йg�B�+3����N�	��	u�g�Q�0��d���A6o�W��XXlxVHYEB     705     250�G���X�7�0���1
�ݹ�vB�J��`����E�ec�ڄ��aH٢�+0���C�˂�fQ�
	4E��~���+|�]�ߋ ŵ�ث���y]�G�/���Cb�0��B�m��r���D��V]h��fcl�B�'NK��I����n�-��f�m���W������de�4���jw4y<d�u[���T,<����_C�VW�q�%hf? <J@��T�Zx ��SX�Qn%k]Մ��[�����R�ܦ��c�������w�>�]�M?��L��p^˴��;��e�0���$2+y�5J�C�z��%_+o�P��ȧ���V�k�TI7�r��S���s+��Cw!�"�["��-���}�����;;*��1OH=�TW�����6��,�S�)LjI=A�\ȝ�4����4�:���������F�QRt�뮂���8��p����۝�5h�By{A���̑�9�`}D���xpƴ�㎩+��J�ު"����>�4>� �ܮ���M����Y��N5��K��ޭ{��cfƝ��qEK���7����ǭ݈��e
��Q�C�	�