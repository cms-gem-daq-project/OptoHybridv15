XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"n��"\�,8�n�v�Dj3�����?��De�׺��1����'$*K��L{\r��P
�X���w�+��ԍq��'�¸J� d�}H�T��GIE�;_�"�<�~�8���J�-�R��Yʩ)R�SK�4O�x[�5|{���	w�������VDt0�6�2^x��� Xp}��֖~yj�$�3�=�݇��N^�W�$󙯱�"V��>�*�q�{h��g?,��{�	��+I
fJ"R��t|L�Q���wS}�%b4�`���C��|��~ջw����ѝ��>[���N/$��J��Y��r>@��l8B����e�ů��m��L���Z�/0:^�>j!O@�j�$��_���u5n���
��7q^��Y�[�܃�7��� j��3~�
^|�٭6�X{Y�@�GG/XLh� �|9x�o)��زƧ:u��=nŗ�1��-�hY�m߲�twi�xSҧ��r-���Gk13�i��Zm���Bl9��Ȧ��
s�OTCeקa���h(<��a��c���<�A���x�Z>A+
|/��y��q�X�{^2�8e���-��r�־��q�����a1�T(TE,f۝ ~�j�SƲ)|�(�n�	�t�`������g
��a�)� �j��̏D���=�=��w�P�v�.=wd̈�ICC&t���%��G�M;r�龡X����;r��#��O�sH �꩝�*n�Ծ�-6s?2����<��I`��u��j�O��k����K�"�2����8$�K�XlxVHYEB    1902     7301<X$W��.[��S$v�nK61��.=��d�>..0'�5���L.	����֮Br�����~ů�픝��]�b��g��S��;��9h�+�v8m�HhtN�I%l��ګ��W���zE�#: 4���&�A�3�~X����٨�s ��(_��R7��k���8����9�t#�3
���ȟN6?��&�;�����]�|�$\�� i���@	��t��r�}\��e��7�f/#��d���K2	��i�;̫��4�>/�Ym��uytf6�>��Ŋ��IeHZK��X�/�a��.�B��f�����l�����g���M�ae�T��?�t09ar%.k�+m��#:���~�'0�}�>y��q���_��Au=��H1|�&|d �WI�v�V�)�i�,
�u�`��(X�dU�՝�g8vZѤ�]8��_�{���b��C�	o�v G����	,ݝ(�������!D� ��Cu�~�/	�DIӊ0~l���A����ڬmg��F���e#��i�zGVM�0� �L* �����̅�}S��=8��d L�)d��#ի3����@��<��8s!���[e��4 Sq��1e�[���W�}^b�6�$P�3!Y|��f/w�t�8n�`�]��DQ�C����NK���>��S"�;�Y���)��y����ڇ�p�q���O� � <�;�m�9+���-C{42d��J?���=a��h��\b�_��D���w��PT�8r �����}���2�������@o5����[�|
�B�~�F:0�G%c��i[m�R&�'����鹋1S���:*��d-��������2��or�F����5r��/�?$�;���HͣR<��r���uU�!D�& ��I��b����6��XNӅ+�1�m9�M%J����q#��E>B���M�ˌ8j(��} ��yf���5�@��=l��jD4����j�0���
��V�8r�\��O.�1Q!`7�u��bl�ޕ��I�Ǥ~�E΂Ԇ	j�5
��f��(�%�#+Roɶ~��-��Rt��Z`�~Aأ_���>F�v���쌣�{�8Խ��M.�
V{Z�Ѧm�T�b�A:�-�DaV��0��"&��a�B@;�rF�F%+�=�!�����6�2��@�N#$/Zr�l9����>>�[��M:a��b-��Z�_w�pүL�&4ھ���WY���^�?8�@)�[44��� �	��]2��2��8�1�fi?�����3�s^!�pF^w����%�^*�|.��HOh����nh���u~���MbwC���B�Ƽ|�o.x��&��S�eQ��
�o�17nN��!�J�f�V�K:U2._�cc��;�N;~u�:u��}$$�� �s�'4���W˵s�J��>���G������p��Cd�ɻ�)"����}R��&�N��FI�4{B�|����Ϧ��e��$ɞy��,\�Ƒ��v3�y��ν>;2�E�幄�{>�nDؾ�[�1R��G��f�n��6��ܝ��i=S��2h�1sPB�&ʐ����*�X���x �I�Ȳز�yg��� �h�A2�M3q�z�x�wb'F&f[%2�a=��O�~�j�x/��BZ��̑��f�����g�p&C����l���b�еѺ���4U�2��6�R����.��)�k�v�K�;���6�t�f�C�=�l.��1��"_�)2���^%�Q&<��V�xL��ٰ���$K$�/,.�%~����0�U����p����7� i��^w�շ��|bWY�