XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|����FTw��P	ND4N������6������b��pt��thI��֯%#���J��A�ې���g�B����Ͳd?���L�3�o$�wǯ�����4�V#��M�DH�l\4�H�'~��Z�W��"q��rá��.��<�f��>����MH�Ի\?������3[�[����)}�A�mrݪ��S��T��j�����n�M���x��ӳ�PR�����@�"�%�s����	�� ��6�'���.JUR}t�l�\�fW�1̀+gq3��j�~'���x�Vg���8��{^�Ⱥ�[��1�A�`nl����IJF�$xl�wAź�Y�P�̓��}_�P'!XQ�!A�o\��P����L��7f)Do3�3���q�ތ����(��|\͙���);���n�j��6_oY��?i�m:�K[�$F��Ѻg!v9�x�#;��N��y2�u��?��q����ć&qV��N	LB�Z�A��3�O2��bW�B��nO� v,s_��d*[*�\��D��i�#�~��;	�ee�������#\N��F����x����.� ��K-�'35\4��S)����_�Ye��]��jF�E�vF��Hd.��篃��='ߤ��@�sb�W�2b�4�WJ�xPE����S���X�P�tX��;���F��Ul_+���5G���`��P�1��ͥ�I�HfI
C������3�Af��Y�|�2��9�n�5��PZ��|��v��B��F�_��k�~z��#���Pݿ�-.�_XlxVHYEB     7b8     2a0u���!X���&��sv�����v�i���~#��	`ȁW�4�_~;@0S���!�J��Iv'�o$�z�[�
w�Y��Tڗ+m��-��ܶ��/a�0��d��7������e��@ FV�=Bn_e�v���M�*����Fm����Nu���_q%I��℗^n�Ȉ�&��!���߰k��?/PV�|�Ӄ�� �s	� Ő�L����j��*�hP���$��xZrE�
�0�m`g��L#�؞x�"ISw��O���\n�+>�����(���$ d�mq"�v�#l�1��������)aY,��A�9K��?'xV���]�@5���Պp՜o�o�������7������,%�g?��E�ux�B1�oY膬�r���ءo�J��;LJ�$��Ś�ѾLHl�m��}2�`{
r���[WAy�:0#]�Z&F��'��Q�Tu^�Q�%�Aa���[���!�p�º%0��K�����h��r�'"Oo���ѕ��	���x��<�ʎT����-�r����z<���� �����eJ�䐰T���cY��"j�&g>h���m�h�����\q�Ǻ�X�0�E�5E��&H�d|�G&�y ���e[+���u���zP'� MG6+�5���JC�1� Czo��q��