XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ź��݀�*V;&|*>���d'�Qvr������M��vr�D��/\�rD�b��.Xށ���̓�^&bӦ:�Ք�`�e���+[V=��$���_)H���	w-ᾁ�9*�E�g�P嘆1�S�z� �yUL��B8�^ y�?��I�r�^FF�~����{���"7r��ԇ��+u[�\�����Np�
ׁ|�.gN��s�s9����x�3�B�?��Q�բ8��bL�$���T��pŗ-�,���%X�q��)��,]�,�Q1������Yyn���g�a�PV�OÚ]���4tl�}^hV�3M�Յ�g]�V��>V�o���nKK���
��Z�Zߎ$N�Z��-eC�a�����\��p ̧hļ��f*��ƌg#�Hh��	�2	n��F)�Y��0(F��Oڰt3�UBʺ�'5��$�4�%e�̅.�'�p��5�A6̙���B�v��R�5`H�؝'Eo7�l��E��(]ڗ�J��i��,'����6���_�N9R =j�$��	��''+�a�GZv��%��H�FX���o�&�`+G���e�9�T���_�������l�W�&��a�z0� d�
�%�'߂�bpo��q��C+���{��L�|�w)睹�n��9p��ecF����ȶ4��tVv$۱/¹�y%
º��O��j�n�m�tT�~�3,�+3�!��@jM�������M߶<�%9��rpJ�i��ޕ�)0.��f��{f+��K3]�zXlxVHYEB    7783     c00���.�� 8�*���c�SݢX�\�3��E�� �(]�*k���j6��I��7 -��U�	{�NM2��c/���`�j��3z]Z�=�ٸ��=F�0�Q����o��7UG�;�Zdk����6&�r�y�[ˆ�&)37�hU���rdmk��Z4�ӋѤ�!��qA��mʪ�S4L">;Re5�{W�&��耹B)}���V��mNR�$��&,��C�<X�����^�L�8�`7T4�_DNx=a���Ǖ%1d�C(��6cQ��E���_.�j4٪�4`8��ʫ��1�p�Ⱥ�U���Iv��h��5�l���V\R3�������u�CVA�v6���K��P�+cBOț�2o�����n���.��qP$Y���B�X���U�����4��ֳ�i&˹0�)���:N�oh^Q�~?"��҈��m�w�N�/4��`�ߍ�e|׹�'���]�v��JI1���8�8p[�fA3ey��d��nK�4j��������ޑ�>�q$�W��+���5���k�Ҿ�a��f#l7��d��[g��6�}���,�J�<J�fA.�n4��Ro���2�Ϸ
��{v�/�;�	"ٚ���nf`V�E81���I+j%{ƣ�f�ck�Đ�F-ɮ1ӯ�A��̖G�����r���B�j������d��\!��H|��@1{G	X����!]��A�ij�'u�t�E.z3\)���k~�T� k�pZKs2�5�וtz��-��Uu�E�7��L�(��8�������F����(��L��km'=\� �i��&e-e��>1�P�.�7��{�:k.c��=�N�Q/0����L�M��NK|�ԭ�#&�c�F�,��AU����K%2��iQ�*���R��S��#�Q����2����S71��4d�JQP�eu��BW�]��0(�K���3mfH2��*tĻ�/ޟ�?4
@�v��#�i��Pz`�#����-��W��{DdEE�aMy��"�Y�ѻ(絥Ũ�(�#�$}b"a��ބ|���F�J�ѥ���~�F2�,��)x����o~��<HNp�+�\�~2Gtc�U�5�7v!�&�!�,Չ�1R���W� ��2�R��̙�+����M2hijRxQd`�6�-H$��]{�#7�9��&��nH����(�d��]��:ȔS�f�,f斳��]�����{�n�HE �"�����%R���.��_�5͞�0�2�n���g�y�9����x�͏(��uʘb	s�u ��|���5�D�ܺ�z˄�h7�4Ew���r��d��<�w.!-�_MnxM�_d�\IWIB�����z��@n1	Y�Q;�Ӥ����w�P;�
C���҉�T`Q�:�����G={Hd^�����vu��z	p`�B���\2�� ����n�+��� ��W%IԶmn���>c`GZt�j�
aB��ᶕ����^�S�Zv��zΝ}�]�TZx��zjU���|��S"[�u|ů�>~+�j��n��n
�y耂oB��Z��Poz֠�#qt�Mz�8|����������{M,�	��s���Ah��ng��@��&��T�	����c=��x���$�;���h�v�K�	s���Ub� a���RX���A�@������J;�W�-��;bk�7��^3c�&�	�̒SG�y�]��vc��5��Ue֥�c.����&:ޟ�OA�<|���<_ ��ѽ^~�D�F���o`�n�RS�^�I��gP�q���^g7/��$��V�X�n�e�I�4q�W���Bָ������jrC��F�$v})�6=@y.l�Ց�ó0@D����q��³K�;�k@	W�F�+��L�CKݵ�E��]�и��K������D!F�㌉G��:U��flI�&&o%�$���i�q,�2�<��[�ȋQRFl��+��=�|�e���&��h��JC�,Uo����#�a��S�owB��ؠ�
�*x"Bx	Ո,�R1���#���|��6&_SuT�M�A�T����#��%���&~�S��˗f�,��el�L X�=�|ȵ
[ٙ��ڛd
��P��'��5���S�T+�^w�~��1���gȑy3[��XX�r�����0�K$<�a����'�����gd�o6�t*��ܕ��i?`�"�?a�O17/T ������y"J���ܞ�]�׷��q�/�n�qK��~Ԁ^�5��h�Fj��g����ڜa���˯q�KQR|�85� ������r�;s�3��֩)�#wv�X~v`2灯�44?�\��0������g�?l�Ij���M�/���0L�U�x���1���t�2= ~�O�:�L�^��uQ�շp3��2̑Ծ$D{�+n4Y�� ��n%3���=Q˯{�]�����/�?&#��v���6�t�%�����֎�Kp�b)�a:	�C�H�\��Ǥ��ۆ#� ���dj[H��}:���"?�8���y��/���A���^�I��-�<��~=I-�,�eL0��HA)��fNC�@��L��*��7���J���+��S]�|��}ּ��a��]d}r��䖔�\��Ƅ�Ň�\�0;��d��$ ص[���J��D{!���$����HF���׌��+�)����0��| 3+nD
�6��}@_h\K��������%����8Ѧ���1�x�wN�R�S�m%;�8��wڊS,%��=���B�P����(�c&�s/�)�M�UR��E��lF�F�l���Xd6B̻��B]���|��FlWop�t}��Sd��S�I`aw��L4���
���ZR�$�)���9�4qK�)��`���ƾlNa�rF�b�� ��>D^.�	d������b����x�cWGc��6�-�c�����.6���;��+�D���[� ��
�#N׏�qЬք�z���d��"HFF< R�ub!���|��M3����\������m��.����
��c0�|��>3hoeb\����1n �xer2��l��-