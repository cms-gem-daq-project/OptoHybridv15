XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q��C�9D�6��[@�}�>�L�1S�iFD=1�yy�R����_=hS��]�4���x�.��U�I01���c�Ȓ����=*��K���ih:)��7!�sB��ҍ����Y8�>Q[`��l�屌,��z�����K��b���Kd��U�7��btS�e�{N1mo��R0�&pL��ХxU�cYiNp��b�kF"��6?�Q�J��*3(	���)]K���H���{��g��7|)�~7R4��}���2L��]˹"��3���K�8*Ov^IўX�h��V��|�3w�y�~~�ֽ��������4-���8ݚOБ�����&�$6)�{Na�*Ë���>1��2�y�fx$���C��R[����ߏg3�z��[���4�� խ�']�
C���?��?~�C�m� 4�p�ln�Yr��":����>�\�>-�e��1?��y�d��1��Y���T�����;�e�S�k?ya7g�B;��@V�}���~�-�i&h/TG0���#ש�������wKy�'q8��h_$�$H��uH��y���M�ǚ�ہ���}�hT�7�N��!j}}Ue{�gC���y-��A�,�Y�.@!���I]�n�ݷbg
Es��|�~,��*�X5�8�(W�8��>͊BS�l��
�"T�ƐgC��|���.���3W䀶Eq�'ی�a���fs�@���;�1�`�I��ۚ�a�6��T�b���k������k���n!�VXlxVHYEB    34c8     730�	 �����ʶ��f��,�~����>� �g�n�����~ik[�
��C�H�Qc��`ɬ�d��� 9ظ30N��M��J%˒^?����ݵ��sd`�&��|��K���������Q��Cؘ_��5�<���m����1�eG6D�	#�w�9p��0I�J:���ė�"g�w�Q��̋B�瑣�FKև�r���X���xۍ����M���!J�y�ݴSm�W��wR��0R6��2I =^��8���W�Ȃ�)\zyמ���������49&j=,��)�<P���ҵ�Mѐ	=�q�bԑ�zE��V�#��Z�\G�M����6�-J,'�7����	�������Y���^���м@�S�A��N���:�����l<���łcg�#1��h%�kil�^�V��"{��`V�������{�J0I�/� �w2�΋�$|�M��᪮&�|�
D�
����w7�D^���KD�?�q�1[����܌W�栤�1��H}aG�h�A�)F�?1���O�`|ڻʫ�$�*&����g�����i�"�|�P[�t������þT͵��`�bA�[=wE�%��L\�������XӼ$�o�/"�a�08�I���d�\�<����\�mj��~.e?�P��mַ��d����>)*8_j��A[d��g�(ef(������P+J�-5�p�N���9�Bt����o��:�.���%�"/uJ5�c����2yO$���b�W\�,�	=`F-��G�j�o{���Юš�"�L��_6���1yd �t{�<$O���$����2� ���j�r�b:�:���T8$� ��-ٓ���/�����ya6�����Gl�Oj�-���%J�d8�Ŵnۍ������O��ӿvHcW辕-�f��
����5�q��r�8�'�����H�@�z)� �+��#a���3匹T�Dp��D����Y���J(�m�l�aMek��e6�Ӽ�W'�X_2h_����OxI	�b�^`o��_��q�`�#>$T���b+�	�dA,b�T��'��.��%U�bι|�"�s�򹡣T8br$G^����M��hWa��T}C��<�j�ʚ��.��i�zs�'���Ǚ�ǋ36��TckNuas��K�F��~��#��׵�E��GȈ{B>��k���Mg��'�V<�XpbO�&�;��66����[$a���T�ꤜ���/�Z(-��WO����f,��3s��H1p$}lZt:�.�G�Yb�	�����mEəG
⿤@:y��NB��8Kh]�hZ�(\�q~�P��}0	E(�Fk�ʸ��Ju�J7�́�S�3̙���+�ƕ�l�U �<z��d���;�'RE�bJD���%���h%$e��I������B��b9cS`N���1�̮��D4�{y���	p�A���Ŀ{����C		��T&����]HfI~j�۩@⳨h�|�i�ECvdP{`:�e���pfĉ��kD�{/Hl�g>ɭ"%@��9dk��V��U<�X��g�q'F��\�?���>�}�f}D�bA�+��~kT���ڀ���Z�Fs�6��?�C��&BJ�ol^i�o4�W\*��m2v	�=����D�͛�F ��bA�6�~� `�ÙB?,��\�O#e5����u��`-�����#��֋s t3�\��F�^�w/kG��+�L���=�=���Dh�)����瀷�M(u�U�!�E&����f�΢�p`��8�<EW�\K8Uī�;(��������·pȲ��<��	e���