XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����q[�������pi��
M��.F�+�gS	����Z�3�|I�ۏpz��x�>@٧�}[� ���a�qb�c�!FT�<�7${/�LqG�+�KY ��|BMI�K1i����ed��pHK���4¢�%��G9�cWD���r:3��)�?���{�;���,b����}����*�e�9�R,�p��䟺� Z�"?s���SO�W�� �O��pQ�Wy��`�{p�����:��,w���W��<G��p}�����h�@A�n�%�si$m1���]��de�	��$.f�k�n��[L�5��;�� /z��i��ʼS
��̸dg���֟�%I³�eP�C	WxrҞV}����z��@%-��~3��Ml)�(�l>�!c���T�'�ʗ��ї)���E�^�%Q�A8��|z��z3I4���u.��mKM�4Э'd�(y�Oź�46�1��8��1�F��>���d
f�流��3w#Q�8jW,'�P���#JJ���l���\ �Oo~��,>k��uE} ���"Y۝��l|g<h�g�ꪔ�i�)���<
:H�0wGF��c?��HfxS��j�*N�g1ojۤ�mB��3K7c��o�i���S���c��@�3�T-����|׆@���Ĭ�A�����6�t�?��*:�y<<���ą��V��(�����dUY��2L�&V��1/���!���&�)��~l�Mi2:�����%�NNϼRm���M(P��Z�_��XlxVHYEB     ab5     420gX�24p�`���Խ��{j�߈1���ǃ������88�j��#�%*� �4��D k���mj�1H�?*�lp��hZI܂pQ��_:����9sG����9.K=��]�[7�Nw�-D�|�w�;mn�ZR�3�&�G�ޝK�=ɇ���-@D+0U�1����7.�D^�픧�_� _�R"�E7���� ��Ҩk�� 1;G:j�h�A�_����;r�p�A��2*]����x��&�V2\��rs��y6qm/�y?�1���� b.��I�,l�.>'��1;lAVX͈$�sh��ƺ�g��;�l��p%<�="_k�b�PD��e3�����pw̪k$¤dyA�Qk ���EC��e4�(���y3��z��c+=�.{f�+T;ڃן����g���F���/|=�*�|\��z�3ڦ�0��qx{���2���*�����!kn2�s���wdV��1�^J9o�	U��^·S$��ټ |@[	�
�*��I;��E����g�&#���3�:�u�^�V����wM=V����%SH��ikľa�`��� �[��c�����HX8���p]1�
�3��u��%��$=����p/9�T��^�ve�܅�e��D����R��*o��/l)� 1?�x�I��M�L��:7quؔ9#����(�{��'"űg�ӯa2`L{�!JG���$W�5����ɾ� l��!��>(sOe
U����A�Z0��;�PKJd˕�q��6�(9ZW�>��t@��<�z�4)���u6>�|�~Z�0P�ٱՂ��  ��8;ɟ��-���@�Yy���d�l���}5��?��Xe��W�x��95��9>��Lat2��yN�ڔ؅���f�mv��֜l�(�%rߺ�xv��ȶ�m����Zy�5��a\�m��2�SD{��K���Tn@p3����D�}���`)>ڿ�VƷw���=�m���Fw�w�u԰<��0:��{��Qߌ���J���#�u�p�\�K�������iNl