XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Jt�-5�����<�r-�f���Т�$�u�?�z�4�h�Q����i���{��I�eѭ�#dq9W�n�����[�>Y��E��zH��0������4���K�)�A"\Ƀ:y�t�nȴ<�B�K��>$�!Z�i� �]�k�����/���KqM���Cʽ����;��ǈʤ�N�HAO�~�\�a��n�hD�/)�j�//N�Y�#Dɂc|����'���M(������jF�J44���R{�;oe�M0a������C��8.�U�uχ�7����f��0����1oš����V��D�s$]& [μ� �O�1I�xc��bL$�	�;( p���|ވ���t��H~�AEB�a����,L�벊f���I��r3�N������,-0��[�Z�k��������Dj'Erl ����Òs~�L��'��� >�,�of �Kv�i@�{��'O�#"�le�E�K�÷r*��sR2��a������T�\���K���:	�7V|�F�5��J3ٕ+T��io�������ɾl)0��G��N��
uj8�h����<��?��H�[��@������R�݁�� WA���q�jJj�n�� B�y8��n�ʔ�R��L��m}cno]kے�o�%�{T���܋&Z7����c���w�l&y#�	�[��f�І��jk��$�$߆ ������:���<#"	a�H��ǊRT�b�.�hrq�g�a��B�XlxVHYEB    500d     be0
L�'�(z�s��eB?�E�F�lQ
.��4��g[:[�K�4h�(��b=�;>�O�X�m�;���4���T~y0#Y'	�X������P�ҁ��2C�x�b�7AG�����M��5�������v�'��3=}�,$0ɟ�:�j�]h��yF�K�z������w�%����_�>%c�#�N*6�>&��.Iƍ�gk�m���,>2zs��5��;��(�hw�el�,zn�z�ߏ�����@*xm�ۮ/UZ>�����xu�D�@qĩK ��(���0p�[���)�����	�w�r/�dR�5]�%}�����@I�0�`>�^��A�;�n��V�RG�`�o+��<�x7�Rd�j��MN�~�,K4"΁�����}A��=Us�a�wg!�	:�Fih&����e�!]'V��F�ɼv���%Ò�TJ�>�P�I(uWa�>���ښ6�lSD1��4�qW��TB�#�k75ɱ�U��?$[ �5�|�
j��F_��m���B�`��J^N���q7��C�ӑ�V9����m1�УpY�7��b45x6���W��>��q�1�ECh�'�०�-0�Z�}�'45ե�V�>C���A^��|�$䫣U�q�f�*k����&&˶�(a�B�T��5��S�:%�%��׾d����T�S��u7��0��<�����d��F�zS&?�Ǵߟ��8�jݡ�w�{z:r퍦pu�x~8��B��S�����%2�������o�j����E�������_��d���x6:��{�"��>t�i�����b��G5�=RE���Q�55�` ���FX�d�D�g2q� 7=010O��'�MO����B�
��Kt��A6J�-p�f"ud ��lMq�)j�A��x6��F[�)8��5mC�Fͺ�mG򠼲�cA��7M�%�`^T���Q��2����1z�)y>ndӼD�E�~uZ�����c�e:�~�]�9���Sh9�x H�)����"W�Xw�=x���y���I�j��i9��Q��_�p����^���Z�^��K�n�a`��3��M;��x�l��ۀ���]ō�%E�#���ȺL�p����2>�ٺ4�/q��"�ZKP��!�3
�gH3V�A��r}�.�;���*�6����&��v
�XHqeA�8�g|e�y�qc��k��7c�V)�>ߠ�z�,O���2��all:�He��EM�b�o�6j[�3]��	�ґ]��u��w�^�0i6
�:m�1۶I�s �t/aAt$V��/�C�-��}i,V���L{��-M����SٳP+v�	��Smg&k��.N\��Ҁ�G_�3�� �~��pe��Zj8�-�,l�Em�w$��3�B�� �N^8���E`#�ȑe`��Lx�yv��c�3��+��w*),tɹ�;T�C�;L\�榻�:��K�b�N;�-S�C�vg��� �H��Arw���N�p���J,������s������zS���)����ߛѾ��.+��^�S���[b�[�6Q:҇~�h�?Zp�����{&4W'T�2v�M���z��Z֯�|nί� #Rk��.E9�T!���O�V�2���y4	z�V�|�2Q,+���v�MƱC�W{ĭ�z!\F�q/���^�y@�ן�ZE��mh��vS���{�#{�h��V�̡�s��2��h�!ʇ	n0J��7��)��J�an�'5�u�nX!y�I��% �rQ.���up�����
�NJa�J'�
0"��t�sӈ�*f�x��\��5d� �ɭ�-V�惦�g����{?��l�]F���7�U�� /j�0NpuȢ���e�U�>FO@���x?1 �������h�1��8�f^�����N��EU̺���ĥë�D}G���ݹ�U�e���Ӭ�{��qR�'�=E:�s�8� �����k`�z{`	>_�m[����p��5�l�Ȉ)�3�&���ʤ�������%�H�J��7b�c��YN��T]C��tQO^�h��h;���r{5�r���T���|�O0r�0��1�޵��dt�V �I���۽ύ��B��P�)���0y(@��+�Q�&)�0�ظε��L��3�#:R]�b�G�Y6|\
�Tn�Zn�A����s���
�?�L��-���ޫ�YA�12�Úw�Z¯'�W����,^]�޼�"GgWn)5vY�'({b��)�#>u���Y�M���u
�ᙵ^}J�Rn�,h]����l$�3iӲ) �*:n=�M���وru_ڸr�%o�����c��wI����]w	�0 �m�`����p
��@k�D����"�0�]���v��H�3���y�C$ǁ�ρl-���/X��1�U��$3��{%��sH��K�Ug�~�@ij0^�\�Kݲۥ�7#f��4ʖ`\VM��7`{��858�
G
Z"�+S����^��G4�en��>_���9���#���{�Ԗ����g-��p>�_��%�!��=y�]���ͮ��O'x�
��CAWdwI���{��"����P�r�����tx�ج���d��[��}c#&��A}.XxjV���ct�B6�E�C�vOm����EmE�=����J�?	���j�X�Qm�~N�`�O��h�˔"��?��duk�'������n0�W�����Q�������zu���##�����/ީ���.��6Vq�E�6����a�����U,���Y���)�`˽~,�>��'���'��Jk%������qS�&����[Q�������`�� �h�WQ�3X�V@���x��� �w�͖����"QD���vW�q�c(�����H���M+ss�w�M~���S��u؃��A��Hɚ���ƎY�\����B���=,�c�j�*���u-KȺ��fP��Ds�D1Q
���~�����cƲN.����L�FȈ�_)��s_��]`��;�[��y/i�*�Y