XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1ֶyo���[�@����@���t(1�i^��d��0_e�(G�fA$��<U.����m���|���h K�N�8ȅ�mq��_L��y�0r���Q��L�0o]o�?-wW�%qM�K�>���K0e��S��Z6��yI�p�A�RbD���4�e{��E�������-�[���e�.\�p�;K�;�X����Wd�ۍ�T�,��_R�W3�{a�\�E\�������^C��������^�$�O9�A��sQ�a�+�����c����W�X�; �v|�+*��f"��H0b�����4�}�����&O�
"���aS�$
�!����m�;]A*� y�c������6n
[���A@��Y1��&�yf����n����9MN39�0@�T�,>l))�:��������e<+g��Kj'����44��9&��d�S�l#��YTJ�;7+��U���
�BL}��Dm�a�	�W�a��@{�9��MO�[�]�3a�^�a�1n�F~	X)�8W�u0��<�Z۷�r��x�H^�n�V@�G�q�m�8.����|{�������� ���j�M-wG��@X���������P�<���4�����{��9����s^�R㻟ڥ�},��KMM���g_)�,$c1t��|EdEٵ�2�	p�e��7D�C���Q�?7�E���Y�Q7�Q�>��|hX���Zs㎬)��M=xx�dF��(��l��U�0�i �|>��'BhD��XlxVHYEB    fa00    1390̀G-;&:�i���Y(��aRqWI��Ro�f�0gr�L��*J�M�7U��4��6�c��+�Q(#Ù�1�	�ޝU+��h>�Ә-�J>u_�w��`���2:�~��|�gx�����A�T�� H�^<.>�+�ff�xZZg2��ݯ�p��X���Y��S�SB��(�E��۝̳)�mx(��"�����~����XH��,���s�͕��?EZC���]RN�xθ٩�̥N���	��8��Z���]]���^;uh�T�٥���H�ʎ���� ~�*�8G�լ���N�d���T�>�lwݼ��d���Ft��/'6�����o3R�Z��L�����:�km�G$��S�bx�2��$���3}Ze �B7ؠԵ�v��rr�˰�����i[�84���*����2V��F^���oJ��e�n�G<\��{1l��ulQ3���g@؝��F� ŵ�@��h����/�J�0��,j��m���r�菫\�b�%"G>���a�Yw��E,��Lv=��\W��"T�S��3��b&�T�Y�	�@�SH��ir'}���fv��,��#�VSV�u�o �Kqz��}�)ǚ�U��R�pg �ܺ�v!���n#�	l{dW���	�m�h�e�,��]�1��Ӟ�#�o1�l5�d��uGbB�r��\� ѪKTZ�kw����O�R��q����]��[���;�b>���l�S�:�I�Df^��v�H�.&7DG*��@�'В�Sࢭ�̡�㰣�yI�[\�H�)�ؗ*�w:�	�,6<���J<���V��p3�.� ��L�;{c��q����l�Ӹ�;��A~p�r��Ok��VVL50�V��(��ٗ�HEK)�*}���Hc�2Ę����2w�`]}���+)���co���_}!���C �Hx3?�-~F:'d�'NY]P��pOޚ��r����6n�9&;x�<F䉧+"���W�I���5UC�n5�=	6�0�A�%,w��r�^=��[��N#�:�2o03�5���Ҙ��rz藩\���؅�f�I�VI
�o�D�d�x��_5�W�@��x���T�G>���V�c'��������ܓ왊j�?��.��ʰg� 5��;ux8Xw��] ����e)n��Ҳ����=����)�RH. ��!0���9Jd�{��@�Otak�۽]L�$cl�Eu�.~3u�8wSp_�^Saɹ#9v��{�>O�������QP6~�D���28$�j��'6�Le}V�[��01m��^�/TO���LL*�1���	�XK���Uc��V)&��u�U]H;k[��?�tX�*��f"f����y@+f���`3gAl��3O�B~J�:��s���u�
�3�6&<'q��y8!e��w�˪�V�o� �P��ex����(N��ԁ-j��L���೮��#T���+��@�H�rx_���F�k^3K��6������o~7A��I�e������N15�^^�����B���k
i� �@�F�e�!�X��T��s�e+~�k=^ew�EU���L�(?� c���0�$�%s�E>r~b��V�ŦozyvERߵ�꒔`�����>������5�� l�ռ�"�#u��T{;vb���R�L�?M}��O�2p(�M�b8��D,<d5J��ߞ���b�c��%�4vC{ ���"u-i����[�1��/AE�Lr���,m�U�e�f�?��2Z���l��z�����R17��:�bs��4�+���n@`��u��*�ָ�7��|1:�K��f��������0�i��$�P�F�
wm���3~����N�)|e��T_Y��_�������o�|ڿ
H��7�)5	��U(,�±�$!p3���bY�`S�|�}q�ne͙b�	��n�A� שּׂh	
��y�emCA�
����+uLiA��{Y�6�#�|����N��7
z�Mn��v��u����FS!�k��
D��O�r�i����d>kC
R���;��%9����%�|#(��r���u���Z{�ihq*=��\ې�r���*�n�ؔ���p.���Ĉ�-���j�S.a���VE�Yw�_�|��E��Q�Qm?j��
bx����4&n��,$*��!�Y}��J�F�q	��SJ}p/�	��rwʛ�et�W����(�ad��&tso�W9n;),̾�QWv�i�Į{>idU5 �=-�cH�
;�1��2]����蔓�� |���@/L��U���3V����ÿ���!_,1�1�&����@�A����M"v$qe��RVS臑m��=R����)U�řt�g9̶����#�_v�3t�>ҢYv���yBD��5ܒ��*�@�����R�A���p3O��>�?�@S@@��	�T�i#ޕkFԀG�"�ƅ�^�@��-������(!#�NCi�xh�^��w,_�k�GR�q˂���]~8�b�X�i�"����H�<�[�ʍ=$�]���.�>�8q����l�2G����I���Ѝ^mc����WQ�l;��R���"jc�!�k�����՚8�U�L܌�W�~��Cj{C�H�N��.�����[H��W��-2,n��T�b�_W�:�����.NK�L���C�������Y�ˣd20"��ĜNc�f���!�#;h�]���<u��b�IOf�S2t��7���m�vW�}������0�$���^�1��j���qTJ^�..��9�:b �߂	���5��� �4��4x5;0-��`LOZ�Z�V��&O��Y��v?N��1˅Pj`�l�RV�O9LK7D��2"�Ն${��R6C񹻐���Q�þ�D�"n�0�g�]
�*Z��E�}���ޟ��Q��[�0N���>���E%�Hl`h��4����ַ7L�b3�g�H�'f�ˍ�dQ,Y��4KQd��9��FY�r�;��Є&=u�6L�7�k��R�lJ����� `hb]������7h�����<n,�b�(�?�y�%�.S>��ˣ���s��^���{�6��b5M?qZ��7�s/��4��F֕8�]zS��Zuy7vYq�/`�E�o�O����7�-�떁�Y"8�Pإ����YF���/9�0>߼=H��t����u[��1��Ł�����K�u΢5@�RP�ƭ�1��KR,�o?�c �����ᖡ����;Kvm�؀�P找؎\U�ĄL_]�}�V)��ǵ]����L�X��!ĩ���tDd�6�ǽ�9Û�":��oлe�@�얔��{�*%H���ZP��eP�=�����_��tK榝�[q�r�IWeWl��f��@g�j.��l�^G���F��B��mB�Kc����1Y#|φ/�e��T���2s�Y�u���1d&��ut��+r��܄
���,4��e�ۂ%qtr�1<�e�/�If�!)'MNTD���	���$�72LX��	�
���t&_[��b��	�Ø�}ܺZTxCp=�^���|�uC���nC���	S�+���;�q���x��4&���sek
��A1�^ ���n�e���ؘ��� Jȸ��5��۶�fZ5z
T�쓝F#Q�cͩ���t ���w�$0IkC7H�Bn����%*�Kk�ص�:���1�D����.����╝�.62�N=I�_H,�C2x@�:�$�ȰX�+�ςi�'h���UW]���
ns<eoքB������cO��%�O����.)�^�-�˫�B���̡�q$����],R���)_q�_����}̫�ܹ�E�F=Ո�SL��d���Z�@���'� ����������&$!Ê1����;�-�\ (8�.5��7�nޑ��W�=�eޚ�5�HIO�F囜�k�*e�����H�%�冹���
턗r��RKg�w0M�u����q�ة��k2�'���i).T�Kf8���X��R�:Q�:�{YLo��٨�Z19~.g�{G�� _�e���8c^��h>cM�D<��V�D�p7ͫ�J��:Y��zT��j���9լ��5!g6��h�Ua��ӛ�_����9:�eT��Ք�U���F�Z�ʦP4�/6��R��J�� �n*ލi4�+�4 ��̐@�?#L�G;xa("|��'ز���C����dV�>�+�C���Q��A"�Lh~��X����`'�6�zQ�+;Ɣ�cZk���G�%(5��h�����C�U�ԏY�<>"ĀA����u��w�'�����1S��)�[HT�u,  .7Zl�Ȧ��"ɾ��;	Eǎ,R��R���8��y��*F����ҏ*cj&���-k�8ĢP�%]���2�7�s���%�����<U6��+�JU�^�O3KYә���T�o�5�՗�o���>=�"��"
�&��[�^�ɼ�2<���Os*�D��G� ���/ˍ��)���J>@[ȟ+��)ܙ��s�~�uL
����:
)D�GO����j��"�9�*`����|>�����v�JǠJ� �	f�������_4Ɲ� �%��|d[I��Ҁ��!z�]c7��Q��Z�����V�`�G��V���?�Y� ĸҮ}s���=@�]U�>�q�G'Gjo}���ٕU�e]t�̞\qg�h(�R�~�`'n�Qʧ��jQ�N�C�/6�u�??t۵�����]���d1D�3�A��':�Ȧ�b>&%��uZ�.+Y���{kF�?�e.y2���R	�y �I���y�6�ׄ1MǪN>��hl"�47�ԠU"�4��E`ִ���S�)����7��0lo^��L���酪~���e�ز��6��F}udY�P�^@o���c�?��#�g�U�u�'��I ��W|�1߄�be�`[���"�	���@�:��u*�o��5х���XN&�!Ĳ��iN[�]XlxVHYEB    1193     3e04�r��v�F���b�������#�nψRl����fѣ�N�П��xW�n;��-@ ������W`�^�$ ��@Su�;ӥ���+�=��Ӹ��mw:�]Q �ۭ6����v��i5��A���-���`Q�u.��Zh�Y!�g��4��LX����udQ�M��H���6hN����-��p��0sJ)��Gr)�8�
Yye�"�(}�w��s
BQ�C8�s��KE���6�����8C��oJ"c´����tw�^�u}�
o1��A�c�!7�x�)��Elr7+vW�:�qǊ`�=E�LX�gH�F_*�9"(�YY�ogܼB�y�[E��^H~�;^�$#]��^�w���^�0/0�c�R8���Vq���Ԥ�
5v=�#x_V�M�_9N�q�o?��h�o���ߪ>�8���!Q+�J&���3BH�#��X.3�6��`�+a
s��)x�	��rj�1����0t_�/�~ ���Y�,�f5%q�ȣ�^f�s}23��v�N��|�~=d��T-���l����K���P�RM�}�?���o��<��42�`�A�D���)X���(L��yۤS6*)�4�E�Z,���fymQSr{`����4�l�u���uke�s���9h�X�*�ӳzr a1�~=�j� ��?�W�l]mS9��ٝuM�7�b�Du�ɉNz�@��ɮ����:me1[���(K���VW�!����T�	VD]�H�G7L�4r=1f��Q B��,kD���%�5HVIQZjh]�ro�e�I�j��e�w���T�M*�395�[WU3*+��^𽸔sh5=��N�(�ʢ!Uu�x�$�xT.A?�2�ޡ	�R��w�����G��������"~Q���l��s���g�l�l�U�6�I.�����4����.�/��UW��1���v~���]�8]�=ܫ7��Omt��P]�"4%|�*�~P