XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����SP�q�ɸ �!$�s��X�.ڧ��b��E��%�c�2Βj�R�L�T)��{
��]�І�O9)T��"��<ķ>!��U0T������=Ϟ��c2�:&�4Ң��D8��H,=���L�:C�l�@ �M��?�HK��xza��,�����9�D��ݲG��i[���Zg!����K���.m&����&ֱ��S��?��Y@���O�n�%��37(�O��#&�����q��5�?�s4Ѧμ�)]aB��,�<&<<]Wɻ=����H�)c?�g$=��7� f:�܉'�ɂ�|}��ƫl����z���a�ܜ8�����m3�������#<��c��z�e�r��iޔ���l�?�f��Skl�]�Tg�i���ހ��32LP�V���#�E�l�m�P'r2u;:�o0�
V����1r������|�6tt����J<-�:q���b��\�X�L�M� �fwx�ᏆX�C�
��EB~�y����.{y�� ��bбV�и6��9I0�K���#�3 6���>(������p���+�z4M����M��0׎j�f����u�X�{�f0B�z{��D.*�z�{��h˓s8���<vK�ժn�����\�D_&�B�[�l���,R`Iш�q���u�š��bkM{��+�W�:�:�	��C�*z�'eO�����@@�S���ˌp7�Zj��۪#I��
����s&x=�fT��SMߡ���T���fY0 6�j���Tw(6�<]�^���XlxVHYEB    1d53     7b0�����t��e�[��<~9uo]{�*���V�=[�d(a�i"i�3�J%5��$|���Gg����7���^�\�gs�x�~�<��X�:�v�6L���>�&�cȉ0�2����#�ڊ��6]BJA5�y�d'ǊP��E"!����	�g��p�I�?&��o��hz��K7���SG7U�bƧt���? �	��]�tv�r�̞12'�d��Hc�y��<��B�^� C�q}��η�"`���_�<��x�_ړhw5V����G9x`�����u��Q�dgUH8�Z���gٙ"�����N�,�5H+��Gh��Q_�0�B�Q?6� �
�KR�F~� ٱ���}2o \1��><�/|1�S��w�a�R�lA��3W�7���`7����g��a�?«��5�I��qYc�o7����yz��Ʀ�#��@ T���eb�`� ˲�#�h)���-�Ϲ���u����i4������t`��B���'�7����s_+��t��,%Ov�w5p���)"T5���V-h��깢�����m�*������>�0}�ݫ[�r%d���Q9P ��~�	*��
c&w�Y$�Q�\}V�ɢH�#u ��*4���5�{�e{�/
��M7��Ue�42���m5��.����=���������?���:T�.��of���9X�����.wS�˻��q�5\ӥK1I�'��JM�����-/'v���g�����%w̦V�����jJ�*N��?�D�c�5(����mn�t~��G���(#�,߽ۧ��Uણ��=x;/�f� �8��ڒ%g�Z��+=d)f�,C�D~�{Х�W��X8 �xU5k����U��f�G/Fs?D߷&� ��ɰ�S3ME���i��e��K�����t�ğ�d���+�m�'ۨS�����p*��\o��a3TH����d���F��%T��߼�!82����!f�N���iO�|U�L梏m�k^�%��G?�c/�~9��H��L�sqye�<2	^R$2v-�ާ`�(��Pe3{pzFG5��U��2ڶ��5Mτ�M�G�\V5r�=��s!4�Թ�z.�a�7�P�ϫŸ�R�j�Kc)W�v��b�:x�4x�W� ���^�����M�k-����8<G6���S������e�&�Dz�Y���nD?�-�h�$�X���8��قM��T�g>�����)%��o&a�n��.M_~�	��N���=J�~I��L�Tn�=nt"�)Szү1�	���J���~7(��jB��y���~WI�����U�v��bp	Ě6?v��}��gvd`�`�C�"�%�.��2�gW����f��d�����%|�!�t���qQT���2�L//>X����0�l��&�h��g!�����]�vKEE9W���M�j���@\Œ<"�r]��_^�����Ϩ�7K۵�Ȝ��cyiB��c��j�H2�k֖��'��,���rU�|T-Q(ƎQ��Â���fo[}����hzV��(���}�;W��Nm�:��{j(�k?���疷ڡ� S����4G�f�zm�6�[p/��}鿧}/�&���^��~��'JF	��&���$����=��֮u9Q?h$��f�o"���/�_�����dcLE}sRhR�3}qF��L���a0XRU8c�$�eJ�m%AYl�����y���G��]{B%j�D�u��s�Y�;43 S��;�<�q�§)/���!��ޖ��0�T��4B���I������R�.J��r=�$�.�� A��Y�=Z�eD�����,�fy�k���� TA�U�bٮ��;p0���m�A���ƅA3�?['���Ů��c�i_�5�6���S��9`}MGH�j��k��~lfGB�>��<Sk&�`N&�Nz��B�OD'�W��t