XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M:(�*OO-��=���z��C��oD�����XPU~�l}&ôTG*+�U�� ����.��>��_�Ѐ��/��(��v��"����.3 �hq:ƣ}e$���ʀ�F���uQ�_���C�}4A${����.��q�����;pp��4J]�wW�S��/eP�l���Tb;H���-DӔ�������m��\U;���A�E���(	��2��xdE���i^a <8��Yj.?<�n�7�fc p�g��o��PW����_� �������0a���ΦG6���H��W�id{Ѕ�P����s���|{�u��7 {'�8r�BGG�%q�@St�~C���	3le��X�o�h��m\/T���,�݃[�r����*��.�Ol�O�,��ʦȎ��{������@"���^m	��dXg���u�n�kwA�X	�Wq�S�*[g)��3���f�{}X\��WSU��t͓�_��Y�(���x���?��2�n\8h�Pb�p郐��� ��ƒq��F��F$V������ߦg��ލk���> ��X%���iwH)|���,[�����L�J+p&���F�+�PS�ku�ı������ǡo�7W_H��S�X�@V�5*�B�����>:�� R� X�<�|Q���~�� o"��e[�noŊ�ǥA.���II�N{V���̄.� i���;hx�ʄqY'�}�W�o;O*�2��9[eV�|���nR�(ŭ���=.���*�iXlxVHYEB    1041     4a0Y�+ӂ�"�˚_���':6 �֩J0��p�:�t�0ԫa䭣LoI#gRm�:䗙8���� ���n>GO�+| t��zC@Q������69�l�r�q���^XXM(�e�5:Nk��}k t�:�[$�_�IG��0����}���G�J6i��=ZND�sb�ԯͲ��v����ւ������/=�e�2J�rhՇ��������kZT��rf�.�(�tk@�4�JXw�� �q��Q�i�� �,����G�}���)8D]��k�buQ¨��1������@WZ��*�J����k�+7�_f2y�(f�o��&]	Q?a��!C��6d�Ô� E�����d�Q�I͋��$�Fn��`9�
��<钇 D��夾�ω�a��,҆�ތ���r��A+lzxu��Ŏ�*���*���^��]tX>����� �I�4��"�\�ls@��-��"�4�nd�[�;þ��uq�:����^��'�Bý��xH}o��oڊ��+R >��W�V��62G3���i �2�U�¯El���T5�-+3�y�shf�O�Z�¯~��dW��zb�#�>������N��,>`��H�x��$�C�ެ6J)@><�)4.pף�;���'t��}��$� ����Dj����𶀽��8���˳��}ʘbi2~���zda����t>���?�*�J��*:n  ja'�xk���9pI��CI�~:��d͡t"?Zn1.CY�%��uX��z���7"n����LXq&-����g�h� '�{^�X���f��!�ζ�����ݍ�P|���JW�������yY�5�1=PD���KQ� ���]����A�̧����^wa^�C#�; �Q��}�-7�p�K�"��xC�\��->��ھӾ�r�GG���,��Z�v��}�Aj�&�YZ�q�=�<D�e�<(���l�n�	(��~����xyC˫�af�!�h�ڠ6h�.���.1��/���?(��*�76N��d���,��^�s�ކ��ǀD�Ϯ�D-�5�k<\qk�ÇO�nB��pW�һ�~n�S^�q62�^� W���w\�~<��RG�x:$m�����j��5
�N�ÙIvKjC3�V�;	t�T�x��B!2v܉q��"��f�巔�7��ns�<�T �uv\u}B�:,]��1'l]