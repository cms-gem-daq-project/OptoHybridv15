XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#����4*9���\���(�}f� [�$c�z���*>�mU�HP���,���IGA�ꁅi��Hߋ��!��"U��+���C����I�%��.y}����,/3��Mn�x�~�Qʷ��3؈�Qp�5�?�D�ǿAhݺ�d.��X��Gn(c�
߸C�D���
P���,D��=���}�ﵩ�]�~k1�k7́��K�b�E�K|��^�Ղ�ɲG�aĦ��-6��Ί	���v�Zфٻܿ�+�rc/����[r�G�17�;kmN�d���R��}O�h�+����ͤ� LB����%��vW��~��v���+zl���/ʹ�����������_����&6[��kЛc�<|aJi5)�n��L�-�<�~��q������Xxن�bi;Q���QHO��!����nW�+�D=3,:���~W���b���֜X7$�+B�d�������?Z�7������ �X@��j�(bZ�E3�w[�i<�|T(��a��~�������mQ���Ml]ֻ�Q5���=�"������U���� ���d܎7�4{�HIc׾�ht�q�/�4��.%��#�����R
\�❗�菌��a��bϦp����/�ژ����`�SȈߢ��f�"�*TQ*�.�&�PSn�d��DET��Cac���˥��j�:�j�<����XV���9�N�������!���e�};-��f`Wg�&�@�T�+���p�������`/�,�i����!�m��XlxVHYEB    1585     5b0�_�c�ԓ����=H�NK�~���Ap'd�x9qM]�������2ӒB��|��21#�;��v�%_���G�%6��d���z�5"|����A���& ڹ+�����#�|�)�� c�!Jy6��/����j[��[�(�Ɯ)�B=@a��zo$�![���n;���A>�,=��xhb��:��|�ҁһ�5�~�--dӐUx��l��5\��Ե�7�W����>�K����Tӻ�*��&�1ϑ���L��Aj��.�C]jb倍�i�Tx�:��������}`#����(�K`�EQ�9�_����Z�^mo��{*<x��E���#����
Q���f�KW�l@��p�c�!��\b�vL}�kBu1�+t��Ba,�6�����1�,��&b������ �O9�m�G7����P�H�8/G� �xP�K��CB��ܵ�w�>�������Kh�Y��"e[܀���
- ��I�:�+�	��Tm�&d��Ρ�("���X�_���j�˦&b��=n�d�o�H����������G P��@�[��5$�,��N�x����M���[:�*{f(�r�@�ӳL�Q�1v� r;E��ڒ����RTp����'CU�x�A9��f�@vv����-z�Iok�����%��˶�iz�h�'�{���>�ɕd�� �J�mQ��N�D��0�0ff I�\�j�N:q9�x��F�Q4LĠy[@<AuUV8�3� z2�� �klL�G$�:�a�O��f�]"h2m>��a��Q��c���ӓXc���Il$ڊ�uJRM�w�?Q{Q���)�����W�;ow>����p���ߚ%�DrD����F�+SC�'ŗ�A\	yQT�W.� �2�7`[��(��J}?0 �)���a�2��[�D�1>6>�����k��{�=���3Q�Њ�*��
<��U�|��-OTo���\o���.N85�X&�y�����J�	5��%*��ȟ��'��0��
C���J�<6e��E�p�U�W�gn�Pg�I/B�>T\�l�Q%��%f�����/5m�H���va?�DQ�Ahx�p�gD
;�d�"|��ip�����;%2i���p��(�[0�-;"V��{�%1
���i�v)q���������aW�^�p��H�b�  ���D�Q_��kͽ>�����H���Oj�Ѱ�,i���W�ɲ?v�6�d�M����9g�j��D���h������]9�e��~�p����
�C(�ν�-��cc�,�Z$0
k3���/�Aʄ�
���Լ�xW L�"ƭ_��WD�hb³\˃���}�L�#���>p�[��+����6�di\B<��xCA&a��f_�"%�_eG�(Z)̍z��Ñ�p��{B+�ٳ��n�ܐ�j���)�A s���T���˥V