XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&c�W՘��nZ'���2�:s�9]I�8��Z��J���码��RD@-ťd[,����SQ�J�1��B��t|&
4�u�(9�DSt��+��n��n�έ|t#G�>�c�"�ݪYea�N�Ĵ�	$^�.��<�������û�ݹ'W�:g���jɾ�E��s6vs���ę����9 nn4l��]�[2�ĺ��z)�e�����X��M�W��| ��!�^�_�&�)��n�IjȜY(�	��6�M<�1>�����[�0b�3Ad�Ʈ�B�^앒e�1�:��O���`�qE��#���3�Rd��|Y�X������%�k���T��U+�O��{���@�挽��gq�����`ڟ<�ʕ��q:���9�̬�>�}�%��>�q^��N>9�M�;|V<��l����j�#����p��L�r^�D�r9��򈻊�, B�;�C�og��|9�Pl_B0f�!�׆�2�7��F){��9�?����]Uv�xG�H�Za��icH龷��_�tQ�s������%)a�D��������OS̈́^^S�԰��K��.�L��*�� 4I5��hJ��r��.���U@��Z����z��,X�s#$�=���g��3�nۉ���Sî�{f�����wd��)�yFk���m2�{��+���d��!G\����J%j�'�(c�|��Pі3�����,��]
,ˏ� ��[����3�d����5tb� A��N����*�~�9XlxVHYEB    1cee     780R��;��'*r�,����-K�W�
! Bڶ�4��+ɏ4wm�/j�ձ�e��"xA��2�+�A^|喌?
�5s�8������[(n.�B�O@v�|=I	�v��E�딄�J	�p�IP�ҳќ{���%^�0�Sv�:�L߳�J�ɉ2���PڀَC)ݟ�:�+V����� .��	��t���s���LB�'��A"L���r��	�Ѫ��WzEFg��0a���������	uE����C�_I���i�ъCHo�#�E�)�A�!�{1�Z��cb/Y�`�DI*>��}��!��ݘe�q�v�,G/�}�R/���dg����<�lj�n&�b����'sm�cf���X��r��k(=H��qxx>���y��ऽ���m���ɩ�!�b�݀�A��g�UI��v��$o�-U���)����V!�\�h��x]���u�ƺ�6�)�>R�e��{}�
����<���G�^��G���*��y�!�pȚ�vItd���'X�i�\��A��� q�WuH�s���ke�\K�7�7Nb�dY�[=�qV��
���/���A��4uHU��U��X4�hs�䰞�oM��
���o�)�7�Ψ��~&��t�/H~~�����V�|�9(�T��?J~՜��xq�-C��Z��V��:����Q�\Y��\n��˩矙�>N?�(M�� P
GP��tu<oX�[�X�]�K�]<(�����(Zp��Y�f{Hq�RZ��|�s�t+I�u����Ε4�}F�n*y�|�Uf���s�V=k�Z2���-\��J�VA��l��g�"ݽ��kOL�T����m����X��ʚ���	�aތG��`�����A꣄x�1��ߊo����&e���;�|�Loo}��e��=�;qkdߠsM">5����A������Sa:!֧# iq!���K���^أA��j��*�����5;��d���X�,�~eѻ�92�w�\��:�$+��qU� �ND�w�%-���t����;�|r�ϟ��d
�,����3�H��K��Ŷ��{�Fi���*f1#��y�,jd"�׵�� ����PjP Fk����%u9d���A�.�� r�V�z�b�sE5Xq"$Z��x�]Ҩq[��EF>'���T�A����R�'��;�Ej`���[G���p�^�QDQ��V����<�[�5n{���-R?��U��Wsǵj�j {7�3���Zm0	x�4��R<��1�����F��{�ƒ�� ��ZiK��P޿ +"_휫=ۢ绾��33�L*��]t&}�L��~��;�*e�sA��55s�C�@���u�U��e�|(/NX9���'%�� j�'�/i3��9���16��m~����@U�5�:X��X�����K�Q	SJ}-@�1da'��O���\S����?�4,�D���[���R�u�{�%��K����+�mV���t�b��
�NuE��_GV;?g���m;��5{���M �������^����F���b�E��Y;�wE��^F�lq��$XAw�v�'a`j��	E]�.��^:<\l'�|�v�h�4�i��D<N>7*YZ���3b������1�kt���Z�#\����r*�ܶ�u�Ҹ	-p�S.��wȆ@�ۉ~�o ����Y�ܹ���7�Ca�U����sjk�"j	�+4���5����_4�H�G�(D�A�C~m�1s;U�!{oA��IGFL�y(��4^�^�n�zRP���G@�V���9��;�	�A��@~
��C,4
^�ঙ��cU��OW@T�:UP����6D~�37hZL���]|�;Z�-̪�S]#��L�@jȢ1S�iGa�B?W3O�b