XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G�R�B�V>{r.(0/������n��?��Sۻ����R-x@3�5a�rxT�U+����>�p����k�
��J��ߧļ`�����R����0!A�yё��?���S[��z��U�&����P2�F�Q��Ӽ��h`�/�U�҄�]p�e�*�� ߾��ҀB[���5F &���_�6��%9@�)�59�4�M�fl����q-wFI�K6�ޢ�K�/���(4u���C��Oߛ�Da��Z�A�'��ZA�C�� R�,i�+!_�g���h�E�#��e�0�&F$A���ʣe�&��3/�Կ;�)5�@�y:񞓕H��zt���kE�؁³���矱��u�2����Wb�#o���n�W��>�ZJ�0�y�����AK����K/L����	��N5B�bO����~�]3`C���(�TZN/�h�0P2I�l/�$�*(� )"}LL������b��ȶ�:�$��Bb2_.q�~�:�B��?�Lț�A�U�E�)\a�DGW*�խbNapJvJ�g��x�.�3��<xîf&r^����G� o�ݰ�Q�oP���&ϰ��;��6��(#K�{�N�}a,;)<�8Gn��b�/�����
+�JB�8u��.���_B^�=�����f3�4q���$��W������k���Bs���9��+w0�N�<�O?Ux�}��D|F�њ�Ě{߇���*'+�Xe�/�b���2b�W
���G�p���O�dTN�� I��@gH_^ I�XlxVHYEB    3c92     900���:dv]�L2 pT=��Fe=��8|ePi:Ǒ:7��܊.� ��5|:�h�,��I�P��]v��`�Ů�;�,�q�H ��H7�(' ��H)a̄�!M�k��^�nM7F1zpo�0�ex>V�4�,�1��U$������o��<K�J+�y�ߖ9��Z&��xܜ빡��) S�7���6Ձ�)2`A�$ �E��?(u��d8+c������s�������g���w�W�Y��'�@����{� �^�`���F�4�z��3�v}G���?��d�����& U�v��{��˙�T�7���ZF�@dڻ�6�wW������Po��[��������w�45[���8k֙�xQ[�}�H.��8�.�s gP���[�S��ؚ�	ax��A��;�U~7�̱XA�����5� ��P�F��t.�@�r��e@��ᴰh�f����*E5��V�|�w�_ ��!���~�s�ƫ?!$��%�G���a5�j��k�(Z�Y� ��j���2A/�!!��7@����T�/�J��\'մ)q���;3Lm�*cN�6S�����޷	I��/�/	�qe+�!�;Px�����T����q���|����X`-N;6*���U����h�d����Nĭ��ӭR�)���"����$.��$���+���������2�}��U������r2��E&���Z��IB���%�{I$����̬,�8%�F�P�9"��e
��QA��KH'���@�����D#��IMpp�9;KW/�.�p>�+:����{�/�����Qx�X �����c��*� �R��%ߎ�O����%e,�#|���'R�l|E����������XG�|N����KU`�`~�'=U|1�TMؠ�R�!��W��9'~,A��:8W�?�㙥JぷH�_������/��_��r�|41Z'��Ӗ�g�ZT&��IXE��9������F	�����]��"���8����8]!vcU���ʃ;����Y͒���/�z.f����t�Q��Mpg�g�`�w.JUqrL��e�'E�\M��;�L�p�Db[�����.e��,�F6���XJԧ������x��	�{d݆�����Vۿ����٣^��IW�N�fʷ�?lF���Fy�H�]ǓU��4��:Z����Aꁙ+&.r@!�ß#O�qc|�r�\=r��ο�d����)��`��!����K::A��h���dR��n��)O���M<��V�C�Gk�h�{M�<_B��� ��,��~N�y�`/���~���t�Km�ȷ/ *>n ]�*��d�N��(�"BsKv�%���[�-a���o�0*�h;v�r����g���[�ϫ�e�F��$�18ʎYAv@��wLm�`UL�f���/�8�y�4%R��������y�^vz��!�/� �w�#ǠSi�q����k�f�ӗ/;@ǅǈ����7�f<0'Amh�����վ� r�|ވ�o ��m]q�m):�L��s��Jgah_�����@c=�F�� �K�J%$�{.�z:)�=0Ս�s���NG��(H�h��o�:Puc����hY�$�c,��@ E/x���$��qd�~f"�M">�R����9����hY6;�g�����t��2/�l�<�������WD
Y��"g.6��*c��D��p,a�s�@�ho�Ma�� rޙ.��[O1I]eҸk��ʶ��B�<d��\���4���1�(�U�-Ű� ��n^w�_lU�N��U�����Ֆ�k �P|`�}�Y��_~Ӈ냭q�����JM|����k�vh�Gê�{���� ��G�o\r�w:���w�w�AX8P
>�����	�������-�T2���Mo�ns�Q�Z�xv��c��N!s�>S½���EU�����!3�KB�Q��u�U��جu�)`��a@x\�Ux�c�k��L���D¥�"tP�Q�a���|<�\�cc��Nj.�˅!�y7A^���9�_�vu��������BT�p�4O��"1f�f h��P������8кJ���"�d���눣ce����%���
���t�]��%����y�Ҋ�s�(- bH�xmp��7�����Vo;�*��D0SF�>���n�{�M
��M��Ȓ���*E%��O 򲂿��wK���uvv�0S���������ݷ�О-m��Rf�͉>�)�Q�:}
��E��hd֭�WO ��E/�� .��5�S���