XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ft�AJ��+�	�L���s�N�;"�������W�>��$����/8�I�7����Ra=��9�����/�w�I
S5�r~c��~�)�t�6����`�/�򶌄�;�/�4����ˀ�o��V~���6X�,�_����)Ϋ�U���w؍h[_I̻0�� �ZLeXVa��8UMo��
���h�6��X��#.�������ҽ퐂P�ß���T��v˼E+�����S՘���h$�KC<V��T��Z⾢d��0SmѣDBk��l8ڒj��1 `O$wJ�z>�4������&e7.発��3�܆)�8
�M�+�tfqu��1`�ӧr�D�˘'�Ϩ`§8��x�Q5��+��|�p�S6���7�B���F�<Jp�ա,�M�r�C��"N=������m��~O���\�<����jpg�s�9���G���8
�;�ؼ��_ȩ�����߲��!�N��F�r����_���vs{n�w���
��
{�oNG.h�03b53E�s�&��J����9gY�~�~�_���1�.��y.�|�v,E��XѨ��;[=gL��=��V���C4�e����!`��11�jϥڱ�Ҿz���d/X�Iǀ�������M�0���h�xi���*�[��UW,�b���6Y�Y|�b��B�XR���"�݊��y-~�����q�3�G�^@du�5>w$���",��n}V��vʜ��=1����TZ�wy�%&g�"��0����1Z�4�XlxVHYEB    225f     610Թ�����t�D2���5�"��!��gN��į0I�/���F͗�"L�j�2V҄��S5#8��,�!V�}@�xP��jM��@���(�6��� �>l2[öaN�'���gW��z��R�l��Xh����A��~?q����"2���U���8:6�W������>�>�h�c�
��K�3�A�kx��7�dRک���L�Z�)c|u\QN��/nzq���\�7��SA�f������qE��y7�|���#9���FX�Ub�Ω>����ߺ��6ɵȖx��\��*W̘B�aW����l�N ��k�"�AR]�3f����w�><Ҕ�$�	��<Li�aUZY�H{������D��C�Zq�������������<�x��x��р%�8�~U���D�3����x�Y�P�L��~ �}�'�v��k4��4c�O�;�Ps��J Y��cY��MI�loUo*Hv�P�	��0��Ù�_�3�S��tEh6o|R���RȺ��[�fT�g:H�*rD�嬺��F�hb�N�?�^.���Gde����=��Q�H��@ U>�oA���w�*B�C���3��C�<2���������WՑ�S�ѐ�<N���m��s.��/�E���
 ���4�E��G�~�H�`{���}����^C���R"��$@���&��^�ݰ����Y�i�{�i1Y,�~� �-𠅽����� /��B��(�����!Mt���_��b�!�����7�����[&���VvnI^���d'I:���^Kl�ީ�)�e�X^ ��F�Wms<cr�՝�8eݣ������)x0<w�=c̰xW�c-� �v^'c�}`�o��"dޘ-�b;v���z��d�'$�}�.���)uMzr��g�"`BC���r啰��	be�;���^��
�2�Z��O� oQ�J?�{���	K�3��U��m��<'����Y�97I.�]q�,8����ѧ��<�i��mH#�"+��@6�	�v)HU�k�,/���	���Z�
��_�3{��a߃�%�w��l�Tǆ7�tq(���9:w�N9		�5Y6�K���9E+�P�#dD?��������)�°���-͋V8�5�p��G0V"���u���Hcͼ��{�Õ��_P�%8�	����g%��/-Y��q��`s�Aϩ���J��Sу�RG`�X:jf���&�Y���Z7�TΏ�-	�=B���O�(l�{q�R:Ȓ1�1�*=�-;�$w���
sr�18�Tܟ����:�@LZT�h��]���X�u��k1�z�TqS+�~�Jlp���a�Q�
�Yj3����E�Hz�th�|w���'��2�Z�a�Ukb�����?;�&>����4'ⓟ��B����\�i�>�R���?��O��E���c"���T�:��l����=f5[�1y	� 9�?��w�>�ה!˘���Ҷ��pM�a��i�&I���s�[F�� �g��4��P;g����t�ѥ�?sF�˟�