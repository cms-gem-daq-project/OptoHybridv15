XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����_��=�!�^��S�T_�x��H`����el��Jvkǐ3�g"�����l�6�����$�z��oH�M��[I���M���Gἓ�Td�����=�cs�\hy1/_�i]����eD�	9rUf3��b)��p�:mS̄�^����<X���!����KA�i8���;��'|�e���8K��c���DovF��u�}�7�q�[�_
>��o�9�����0r���,��M��ڍ�6岎R�x^�B���9�+��9-���Jk�����O_��߉J��~�'�l1^����[w;�;�=M ���˰s�	���^+!�ry��˅�~��*zf��7s��� ��p'�]�Q�%��(�TE��d���Q�k�9����SI�����1��� �]��W��iQ�1����E�-l�a���UO�9,o�+ΉRHn}n!�7

P��<t0_�[�|u�»���佦�����/_ٔ�	�-MEC*�Q��$h14�ad�d�07��v��u%,����!�T�z�dl>�t�5N��ʥ�!�1�d��*k�˹�V8���o��8U�\qg#\]2�RA \\�K|��7���#N}���_o��3��%�X �х�Dw⌂~�^�v�
��8����S��$V�}?Ϳ�8����F?�����~�([�wZ{��K�3c���_��۷��ب��Љ��@y��F/�RA`B��4�6�WP�y}�t��ժL�}/������w��*�˕I���$�PXlxVHYEB     ddd     4b0��R��	�ZJ*ϑ��^�\�'2�����������Բ'�S���U6�]�2��&����M�(��4jP�/s#0�3V�
b@Cm�ڵ	����3�F���be�1BV�M��,�.�ۏ��I��j+��%5i�%Ǳ����_6���̬�Uo�؏q�=�������#�T+=3�g�,G�|�9��1��VR�E�E"t���b"�}��9-�Q&��Ȭ�D�<z ��l��n�_�m�na"����0�T��(����G�t0��ٽ��['����v�y��� �MiG-��L�2��( C�5���j#J2����EP7��һ�㦎$��i\~��T:��c�l��6���xA����:B&���pT>7v�RM��[�9:����.��R��%-�����Aصu��s�������$^|�R��7W,SV�;f�gp^��@�V�[N�i�/v�O��Ʊd�X�x�d)*�q����X���w{��!�=��K���dJ�C��&HM���_s�+��kmr�֕&�M���M�9����[�G��;Z�s�	���MQ!��m���;	n�"�Gd|���ZF�������,v#�<m��G�i}0pO�\�J��\,�BN�NtM�҅�+-ԙ��䖳�	m����H���D��s��2�>}��g��o��=F]�H{�55����a��EE	�>��c*�E\�e*(�!����h8�8j�ޔ���� �iO2��ft���#?�S�7<9��Hѡ=gd(Kk0��9D�'JÜ�g��ZH
m_[ړ��ڠ��H8"�D�(%�|�� W�u��sR�M���[�v���k��m�rs��4�r�d�XzW�:`i�mOǤ��5�%��gW�̊
�o!(08V1K�\_��|�^՛[�n_%���u�����	a}����xK
NU]R��)uf*f�s�߇j��w�n�a���Q�G�(���B��7�e[gF{�C���<PA��J|c���U����n��C����H}k,��w��-�k��:ń�*���pb(9���,�&&���#ps��]Iz͸_k���ѻ?e^$��}��@@6j�9�Ͷ�t�x��=HזB�x�����xd�`f%*��u��S�D�r���/�158�� ��̰Z����8�Q��x%�%o�[[)�