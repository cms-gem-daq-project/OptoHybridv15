XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y(�I*����Q(�����l��� =T�{ �ƾV�B����eZ�S	gq����W������� }���/d���"��ZID��!%́>'BA/��e���6���X���Er�?�9E�J�3�^lP��ΐ�2���UqZȻ�n{Ėp�Pt/�����"p���c���{f�?̲�n��c0��Y��e�9�nc���	�4j,Ǖn]r�US�f���P;ĘP^d�I��>�� @Z4�~�塸�*Y��b�e���-�n��w��^Q�󘜾�*�ьq�������vC	&�D�;��1������f��{l"]�x���:��t�@��Ձ�Dm+��c͊�s�ǝ�f�I�@&"��*�!�����G�?B
�s�Â�4��yӕȀ���f~��p5�}t��:�w��mvOI�7p�ԗo��hڭпh7�47yx�?�����2mEY����X����O��2܈�]��M�\��n�Z���O�w���Pw \^�z©������Ӗ� ��HIi8��Y����㗶�|[��v,���<,Ur��U+������@���nJM��h����S�pd�MEc8?��4����+'�΀�Yk�L�)竗�9v�O�p��yM�%7/�BwY��@=�yCy*�T�9*,d3m-<$}�,�³S�l��q�QX{�K27���"ɛ�qV�9���t����E���agU�@��(¤s�;(�^o��d!��8%!�P�o�K���{W_�X�������,XlxVHYEB    1392     550�":
7���l�v�w�򃔎V��&q½+��0��B4��L�wrd	�-m���R�D�I���_�2a�	lA1�X���Yh��%��d_�U*0�܄��8�h�3�r�mN�K1��{���*�&�@k�m�wg ���3�JX�����蚶#��4K�VA���_H�fN`��7�w��+�Zd5�0n0��t�=�Z�c��_S�O�].�R��)�x�ۏ���K�?�}�C�l�l���0�済K�Πl-��l^�U��͢	� xjs5�gl���{{�
�R�骁R�����!��:r�:��b,�:��il$��!��t��I!6����#vq���-�@�e11�e9�o�����ʂr϶�7�?�cs�X��K�}Tݜ�|G�<[2���r��	��y���l�Y/|� Lo���E|�����[
��	�C����`(�L��`U?/Qo�pP�p�x�w� {VL��n��i0@�q��D����V�V&��b,�{f��@{xX�r��Te!jv ����h��+q�9'�Ww@��%��9D�M���V����^S���d�3{��;��~���Ӕh�Hm-���m#�O��|��o�;����V�&��֦�E�>u��
�3�?��8n�3��!eyn�Pǚn��jh�;~_6}{:��J1	_�+[�魱R�F�l1,e�/��T�$i���L��#��\�+6�s�H�>˲R����cä�f�M�I��nr5У1D�Y�_���$�ǲی���e^R��c��>�0&6�Ҩ�1��\̀G;���՝�)Ⱦ�q��DU#����!�1���ݪT�����D8�p�(D�d���ЙY�{R��1�4�P	���F`ܖ^D���Ji��T��跚�Ve�ﭴloɇE}?�̱�о��� ^V���m��zXh&�(qؒK�)E�
��
�6V hj��,h��k�3PP3Ә������kur �{RcU�Q���O߳ȭ��yj�6a.���9S�&,�7w��a� �<��"�f��1�r�U�<."�n��#B38�G�	+u�}�ځq�!���e�?7�-4j�����ţ��[!�5��gM<oO:<C��evd��Ǩ����D��iХ5�L
B��<��@��-툹tr�3U
����!t���	�hF�̝���1�9���ԋ����q�x�?�@����I]���~+�t��ɵ���Z���x!��3.M���ҥ��B�@q%6����/���J�|Ln,_�Z=f�_gH�l�Z"��Q�����f"�;/{9'���J7��}�d��F���o�����El����