XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���eF�A+3��*��JR��s�<x��ϔ����5����_�D>�_1���}I�K|S1ƈ�֧As)Z+��8�ݺq&�_B��q����0d�����������s��)M�T��ٚ��z�*��V��q�'�e�+s��F���`�ۍ��R���Q���q�W�6�5���V��5���W��U'ղ~8B}6�'��g�%>p�Ӭ��
�	o��-0a��k�����Du���X���h�s�Ԏjٌ�2�*C�³L��ۗS��FD�I�]vH�V�c�p&��Y�|d�T��	̣��|> ��X����`=��Di����.��3�T��xB���ɰs�л.b=�A��'�5�/	������6&4q�RR�.�>�M!�����2ƴڞ��g����)n��nlc�>t�V�F�2�2(��H3F���:��)���s��lXk���^b�Bj��ّ����씆�&�~�����ux
���A��������r ���r�����}��%rH��x�s�J�$��6�������Gf�D�UL�ل̓�$���"V��<�d�������ɥ�t �I<H�����R�x!��\�f�@[j�)� ����ͰkD�O��]ݑBQ��@�Ɨ:�A�k8�H�/���א�E	�q�#�vqQ�0�:M�ge���n�p]��m^w��V#[����PΓ�k$�dd�8�Jp9�!���5E)aS�~H\�=�z��Q9(�+=-��vXlxVHYEB    1491     490ϩz�§��OΥe�KՐ����y:5��ꇦ.(Gv�V�a�
^��_�7p���w��b��S�d�6�w�yr�̮�&����lt���� ?�^%�4J��j"C<��ؚ�p��=4�s�Ci�������y>6|�7�@�C'Ǎ��7����G���C�ĭf!�M}�3
>���e�G���q�g~�*�"&bȨ�ġ�(��'�,��ӁG֍�~�L���l���P򝷪��zoafw����{�ކ�kU��[��S���s�d�8��QkZ��C�����ΌbH�U����ϭ����va�K����q\��T�#!�[{p��ë���q~!2f)�s�u;�*)i;#v�)9�}����>D�oa���ٵ.�����pg&Ȋ���x��{���_������0w*��谯���.��I��C'�Sτ����G�)o�dzE��Sa0\-�s�F�2Ɵ&4����r��\,	�a�cŀ.�.w@jV���Ƈ��Q4�6��)��-�߫dc5���CL���Y���hS1��z����Z]N��2�X�uN_�*��@�އ�-9ګ�ʌO�2$�j
��6d@F�Sy�7���cק�B#���@��n����5��
�6.�H�w�ۦ/��9<�!�;/Mz< �K�M��\Ϣ�HJBYV�xD���J[��knG� ��u�F�mavP�xg(�I�E)��c����#���h�<?d�1˴K�m��]��`�)&��_�ފ/y�b�
9V�H/�ͮ8A�^V!�ȉ��%5��l�k�F����1�ۡ�Z��wg�X�ض}I��]�}K\0#�4S%����c
*�Zw�)U�����#�bq9Cj��S���>��X�(M�����oJ�3� �3�~�?ohr�<��\�����>Ƕ�rq�m����p������]�^�`���kِ��*��Ԍ7V���Li���ߚRSW�$�{���-�#�C������cy��tDl��QP-:h�����O�ۚ�������)�����N	����
���5F��-�l�(��|a�n;O|���f^���&BT#����A믙�R¤"b�[,Y�X��Cr	!˙/��(hIv�����<���zB�/D"=�&�SƏQn�x��Q��?�