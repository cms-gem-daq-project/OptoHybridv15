XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�y�����T���0���oAj�������e�U�qq�F���3rz�q/��,*��td�L5��ln��:�.<�O�J �"Ke����mͪ.^�`�2=
 G��u�G�v��י������	�auL*`�%˦��:���h�@�kf�ir���w,�M���?X�N�,���H�j��n�h�����?���P>'j0ߚ�Lؙ80�
��N� �Jh���O.uz����`���[��!��r�2�SYI��r*�)����V��Tnp��١�����h�&dp��9Jr3�/��ϦDQ�?c[�K�k���Uߥ�]��,`�*n吪����=*a��]]0�j�G4�.�Wv���(������_��P�h�74��[�C�L@A���L�t7����g��_�&>vc�;�!��7�n�	e�a�^��D�M ����ѯ���w�; 9j���������ȫ�/'�BK��?3�Έ��]�(�s�Ď�m������%���4�O�f W���7bS��*���.&����b���	���������}rQ�G����9_y)���� �v�;��+�!]�՞AuV*dV�Vơ4�+��"}�w���-�/�V0�L�Ӌ����i�tF]�0G��J�R��}�ơ�l={�?��ETS�6q�^��9",I��@LI�#�� �o?�	͈�W��u�5"���<��݋��gᗁ��+EFw���0�dB���53��7=K[:c�*�uXlxVHYEB    6fc6     c30��y�R��(-�~^�*s��*W�V�WtǙ�z�\��p͙�<�.&��+����$y!��@)B���%�F��,�8�gF�T�6<?~{y�_N��))`�R�sY��H�ByRz�V�4#�)��j Z�Y�.XhĻ)��GYF�L���Y���L�Kl������uW�:���,�[�р$�D���W�)��Q���=4\���Y�!�x�kW�V.h�%NЫs�C�_�O�r��ڽ�:6��[�cn���k�.�~�֚6U��4CRW�W�â��s�r/2�L�_�þUh�-w���F�&/4N]S*�X1P�TU���ѝ���_��Ñ[ah'3ad��%��g��?�K�\I�q�P�,X1S�
�h�L�Y͍�ظ�{��[�����A����OT����з'��<i8^9O��;�/3�&m��z�v]������}��,�.6�\���.�������¸gw��u�j�Co�H��n�!h"�;O���e�\�W�N��� �t*��p@)ڒ8�p�@�`ê�ht׵C$;98��WJֹ^N�S�9^��:�a:�abT�����3F�/�lM��E*]��|�� �F�k�ڭ���W27(+C�z7����[3�z����*f�xo��?�0��sVԥ�;N��w� �H��R�����ɝG⽏�T��tg=ޥv1 ��`���_B����f�<mk�ž�,�7yMd�>^z��@�uW)h$s�	�	���/{n�-�M��_�5�j��&@td��L���=_���:�CôC�����mIf�5sjws�^&�l��M������I�'O�:�Sʞp.�=\ɽO���+��pI�j��φ�t�(�!n�HT����_܃�v�hZ�CT�(׌!��
�vm	_��P6��e�VG_�@]�ї<�O�hli ��!����`xHO~�5S�&S	�g��2����d�+�%[�iP܃`���~�RU[�Lx[) ���N�v�[�f�o�4ռ���y��k-��*�D���Y��ƨ���t���i���iFě~��X':��T�V�'w�?o	Y^�Ѣ��0�_�5ߝ�7���עd5�.Q�H���%ե����An��MO�`|�Ɵ�}��	�ک��ˊ��OE�����$И��u^-.�6��ܩt����5���s?�_5mQm��I4������^]�s�ԭIc�w�*,>�˪�Q��h`Zy��;5M�=T�,Yb>X�ŷxg��=��`=F�q���^
U|��X3坞A廁jg��?5�O
h7�j�ǯ�D�	�,,��X螒S/��VO�hv�{�������)���Q]�n���o���,ۦ"�ꤵ�U���/�%���c��%�Z-Ȇ����R2h�97�W�s��ˡ�(յ'�p�7=cPrN���Q�ágW{�v��B��.]:?�nXf��z;������e�l+�o��
��?��8��)A�z���*�Uc�9_/����fҽ�YJ���^��=?��/���'y��η���: ���ޤI�]���bG��|b����Bۮ`i/D��b���D$G�y��#a�H�����ϻ��t�W�� ��NΏ]Rh��U��煥�$����.ҩN�ۄI���q.����9��:�!���Ľ�8��aFI�D��9l+y�xE�q"��"t�97��C�jR�C�(��D3Ji;,�m �jw��>AO<�P�Gl?�aatZ�G-������:�zŶ.0���Hd�2z�RH��N���H��a��b����bvP���aqz& nf{���<�\ZJM������P�]��J\8ܩ��N��Ec��)�rFYd]9�+,TM�/y�u�8��	Su[5W�Ύr&��;t�3�,�����ALԉP��OYB�/`Dh:��C����㴋�ӏ�WC�JԀaïd��_L�x/L�v- Q����Ȩ�
�{H�g`�� ���p��R~�W%e�m%�ܵ̈́U@�5|����x��[���a|\�	)4�/�A�q��!(���}��4�7=0n#s$�K�-�����8ZѺ����ۚ��g��qM���֐E),s��ƺn{L5#�'��)p�TA��yb�2�ŕ�?��u�a�'�ʕ��+��5:�Mg���)����[Q���㏎qژp#.O�C0�X��sn0 2���PMp��OM��]�$��s�&X�<5�$��?��v���E��}!�h��I�ގ�U����W�At���i������Z�tDy�b�*�0�&���V@g�����Y�S�dٚ��40O�]��P����9�@�l-F��L����P��~5�u�	�Ժ�n�C��ـW@��Y�s�����T�	7S� w���&f�/�uϐ���c6U� ��0��8����T�mm$Z��5���A��5�<\.��l �x���`�(C���R���񟓳C�l����m,�7rd."*�DZ��.w��-��݋�:�_��p(����I��M��:�	��5t�6��U,=X	fH˛`�ITN�jI�$|Oc���a���K���l�T��G@��Ӑ���S���G�0D&6�,U~B�e5���J�{�\����u�Ǫ�g~�Z��lϭ�����J̷<�{K��4����
��)�!���,�<�5h��kF9p��y�7�	)����^V@k|1t�׆R�\1b��uN�T�����֣��������c��E�zTU��� B�MbR�4���#	�F'T�re����)��Y��qCt�-V󷭏PL�Y8�w�ϐE2ذ� 'H^U���.��ǎ�JYN-�$0�� �~�	�f��`��!� ��l�S�s�BՋGR�#'�ə�@�U�ŧ�����(�%}��ȁ�@�o�(Ts,d㐄�c��D������sݟ��Șaؖ���=�*kdg�B��[s ����F���r�}O <�
8��/��)>��Y��h~ܦ@:"d>l(���LL�m�2�K���w��Կ�Q��R��x�0�p�-=��Ls��;�8��C0$oO��B�kYg
F��g