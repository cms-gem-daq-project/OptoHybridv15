XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Sz�&*�(�@��L�A�|u2 ϥC/V��@�^�YM�j�1�`�jY�qD�Ŷ;�x�ϭ_zA$:�l�� l]I-�9Cc�&:P�çE7cy��Ԛ��Q9��⌸Q��hlQ��@�G��F~ĐQ���
�9����`�J�e�[\��I2L����R5�Hߑ�\�9a��5q��{u�)6�����0*�����+�T�r]3�A����%a&�Q�9�f����q3��R���$C@������]]�*%�<χ�1�h�U�/x��V�I ��������Ը˒�(�ZO�$A�k%-�("%�q�^�x֋.�
�b���Z�	K*�p}���F�V�������*Nݟ�ڞMb���W���Rd(����e[J/�����F����[q�=##���GH����qc&#܊t<�8�m{f���1(�8��Ek
۝�/�G�����$%�R�WF~դF��%�C���6^C�6>�ix>��FO+Z�0eĢ0gNt�ذ��@�G(>`��������R�1��Ֆ$�`v��O9."(~u;��}�Z/"�޶;j��	+�����U���o:'pyT2p�6ߊ��(R(bI/�B�r]-���.df���B��:�g���}(w{8"3M`���U� ��9$	�.sm���T�=33�0l{��_ U����]��..�'�����p,�πz�oH"���]�h��I�y�$� �?���o��|���K��΀���?�e8��M�="��]XlxVHYEB    2864     8d0����[�!�ݴI�ʃ�)��F?��u��儓`�*8J�u��Hx��I0ʸ�E�pm�>;$3���F$����ؖ�JР<k�ec>�;���F���a�2�%&���
�w�R�!�z$A�[6'͛I�#��m���#5j5�h���
�c��Q[�u]���z��R��M�����(����឴CWH����&� ���K��2��ae"i��E�l�z�����c���,�ݖǕ��p��u��Yt[t���
���sV�"~T�+�	ߧLgwQwVd]^�TAb�JY��5�YQ������?��⏪^��e��43OxCci�Pʁ@fY����'�L�L���`V�Rv�n4�Au^"t�/b`b�Ӽ��C�1��ՐR�����fz�e��v�P��V=��[ƀM1�D��(}�<7���'ˮl��Z7{�q:~�o��'q��
�J�˟��s~/j�AE�H��]�bdܷ���8H��Eڈ�h�;|֤ݴ[]/}�8�:"`�ȼŭuNjb�do֪��rF��d�B=[V���b��r�-zG΂�4#����R�노�оNz}8�t��C����IC�kLu�N%B�}���jH�d2@x�ҹ�Q�y�k���jr���f�W�^I���Ƴ�8�G�Gp�/��Et�?Y�KI0G�P J+��A����9�w��S��pq&���!q�����,�8o� �"jp�ϖq,�UN���ye*W)E\-���8�|H�L�}�h��P(��\���SQo�<֛=ٷ��%�
�,���z�:CA��YB�\&8J��eͨ���Eg�)J��/�c����Wg��z͙��}�,~�nj�i��W�7,��gx�I���QӢ�����J|��y���ޅmD=�A�%��I&��n�>>��{]{T_ș-n��T��2�TD�'	��V4b������]K莄�%:r��!�$��춶)9�J�8ξR��`�Nj	rk��1�\��W7Z{<��|�xp��=($�V�"ۨ��T)���;$���ඩ#�PH"��i��1g�����Jhi�̶�l�o�Y?�����6��G�����HX���a�+PG�H��U�P��)��<H$��!*XU�ָ͏���ofY��N�l�;�Yp��p��%�l��D>}��"ŽB������$Y�p�D�51�Z�r��lIk����k����-c΃m1 r0��e(���R���"�&�D�����~mU�m.�R{Kޠ=���RTX��C�[����, O��p�zW�~�I[	0/t0��<O?sI�����v1���*�SSu�YKiS�����4�߄F?�}�(���!Fy20/#ۿ����k�m밧���F�{e;ѿ�����'��_�Jt���[�0u�B� �Ј�qiS����>�8ަ�1����!A��v/�+W/F�CS�,'��������W���P8U�MA��~
0a��k�Acȉ?��+�FR����$�q����n�7NK�m�*�ӥ4�`� ���Ï'-�.���Ϩ���uDD�����y��d�Bv�m?�f�sNb�9�=\�u����(�H%�GyZ�_�A��l�L����(��v^��T#�����DZF���}�DT�Tl�"oVTJ9U ��Pq�:Lb�hUL@��`B�܉gw��? �'�B�� �?^�����ؔ�|w�h8bOA� 6�������ЄG�5��a��eC>�d6�o<Df�����G�7�܀UJ�?쟱c�@0�l�A�[5	��]q������E:�W�=���ƽG&%$��<�w��~I�邑=���s���W������J��|�����4V{��>��-����;5ڑ�m��j늓'3�GRר4(�0�B�o�!���S�o \�l�Q�S^@k5���]�H�K�4���45��"��?�FVÉڦی���Y���g]i?j��g���[/G�1�E�M@J��\�#F7��ΰ-��t�c�h�Jy�'Jq@����K���Ii�"���Y9,�����Wc���=M�C
������M���=��)9��f�^bM>��4���㉮~��*4�>u�և%�(@�-6�k���(<�V{Ts��ȯB���@�����MH�#!�7��
N�E��R�7�8P��8�G��+�'�<�J�A���K7�v������\�A��cR���K�����72Z�*p��P��W�*&��i��n�*��3�eC�