XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����q:�F��P��h{60���r��F>G��Y2�
�_����O,������)��겐O����B^	l����iT��!��-�ݯn0���&d �9�����A� ��]�����z�6vd�iP#DC��]CM�H �,6S23v���� ��)�������=�4��s<��W+�:�6�XuV����?�5]�%2���12��r ů>\���" ��s5(�[.eB�KT0�Q���?Zy�\��4�G �PI7p>F����P��2�r����%�s�\��Vu��t, ~����d���_��WZy�H�KA�[Ӊ�(/~�p��9�#�ɮ'�:�.�!�Bӵ��m�&�/!�s�b9�����h��:D�!���/ɻh�_L����@�q�h[��=��vo�*��)DM+�w~���kf+H
鑭��޾\�k��� ���Ckwya��E�~��T���^����&�7��W��M%��Ȗo�fm��M���>��p���I�	$�g��k<a/U)�io��U3(��:���k���������[��^�e���pWĨ�~ğj���Z�EQ<	���/�� ������~'j�
���X|�`3 �=�y��6�:�%��K��$?aO�Z����<Œ���ka|5Hj[�,s�e����c9A�[iC<˵��%�;��ۡqN�V���[�I!�=�Ayh���R �e �)Uz
�)LTP�!�,�{E�>P���_�TXlxVHYEB    3541     ca0��އ��y����ٓ�6f�MbQ�#�.ҹ9�b��d6��V&^|6b���>��н-ڪ�Y`��+ϟ���kR��G��Û��BP�a�:�;���_3ć��FȞ6T��(a�?	Fƃ�:�������GX�1P�f[)�;�q�fg\?E��[��M����Zm��y�d��Eؔ�����Wz�w�,f�%��x:
wVaE�Ѧv�Dn�H�"�G��N�`�Ğ��HC��A�h�<��m6D\A��$��X�QB�
�>s������6E<��,��I(���r��|X)��.��OգZ�X��Ȱ��ڰ�}f!>)�+�U�l�5�
7𡜔��G���Α|�C:�nm�8�@��K1�}%^�nxK>4b�D8E���~j�Z���z�����������v�1Dힽ��3���i��x�uEb\�cb��.Ri��v�0�|ꚉs?<�F�HS���O�f��W=��\[�eZ�~�W�{���]�(C_(��-�92�iu1
���z���+!�(P&�DT�3M�2^���������򓊞�&�6v�q}�ĉ:n] �A&��"[3�
�
�m�3�ˎC`͗����dM���i�����_��W��j�&�M#����ԅ�01�Z�|��Q��(X��XJ�Qz�%��iF=k��x��p�3���,0%&QEYj{t�S��~�����P�G�/���[�4�q���T-��z��il�dS��:T��'��Cw�|R��
�����L�w��v����m��öF6�mJ�K�7�X5�-V
i�����ۤy�RT����v2!ڪ�ў �D;�#0�㔼1\��yJg�<L�}QA�`t�p��l��o6
k���h_�x2~�V7��|#�}��}�M6�tq�/��VM�ʆu�Q��_fnq��v֗�+����}Mtk(G9a��.a`F�֜�ԥE �tE.��Z�Ub~U[Z�#��I���|�x���iЖ�N	Ì������q�(���	�.��%K3���i4wg�Q�V�&V(ci�-�Sg�]Xf��Ĩ?d���+��;�}2�`����5�?N�����l~�hir����>�uE��v-�Ge}����3%⯁�w�;�J;���.��V�]�}�Z����#�tb1�d'̯�=���d����;cޙx�Sc����)��5^E�L�>6�}�6p׮�:�ʮ	�纓�yi�[$��k�;��o���T�΁V2by���%���]|�[�goH�ɆX�,Lt��$��2Z����|�YXt�nC��
�0i@��f�T�J�H���A�籭�cUf/O�a��9X<�1Z�`DS�:�	r������˶��ЌE��B�=o���Ǿ��*gG��<lS�Ǧ�	H;�R"�dx�6��(V�aI��l&(�18V�(o,v����PW��9�˞(5��(�{?�@�w�9��@�tE�����m��83U�]E�[Ɨ�1*����p&��^��FR�Vͺó��y��L��I7Ń�&�2�<He5����"�;{GX��Y�_ļ�I��}����[z6�U�	LH<˹�i0��@�"����F��5WQ��:��e�B�%��J* %U�J )�=�mv�@���u�zR��(7[0S�c#�08�q�Rʴ���b�Z{�錚���^�\�7�V����h���Ƶݢ�6K��w\'j�� �c)�����Q���2M�P�����}��+�Z@�����8��0�;gD�VE
�1�Ҳ���4�إ_�	7��H:���?��w��LG��;T��vs��]���h���F�}��I��~t�X���%���?HAu��J�	�d_����>.ό{��6���,��I"AFk�)���4�����U*[t���'���#C�76��6&���F~�N��3���x<N歾���G�ܤ2E?�!��-	��'����$���"��6��m.�c�'��I��'��/���ޤx����G[�j�'��ĩ�庰N\��@x.v$S�`������N�Y��,��A<l |��3ζ:��_�s���ͨ��D��K��:e�[x��#S�G8�j�� ��	�s|0m�"�}�|�#�*�f��<��I�9�T�AВ\i?�#R��Z���>$�@���ʛ���J�i��k�vc����µ"���c�"D�	�{�4|F�����F�-���:k�ߡc6;j���!f#��C��l�i��38��|]t�l�ȤL9������H���Py���I��ɀ@jD}�Kc�I�/�i��Cr�� %o����	7T�*��Q˃����U8��A���jҪ��}E�E����ޑ���/f�z��5�����U8�m�X!�Yu��%�Q~��7�O�rwA��6�m9��l9j�]��z�j7=�N>f4q�
���\�~�x�kxK_��%"Û,yR����6Y|�;H��T�լ5%OSOc�-����8�{��=�RKpX4�ݣ���'p�V�D�Ǫr�u�t� �>�Z�~y|Ô~����7�W�*���U}[�����)%n�8�	�F5�$��XKd�/�-Q�xm�qj�`�ۓ,��T��Ì�VTh�k\�G�7q����i��=��Z^���?�L�դ}hW�ej�KD�F��g����G_��V������|q��2%��C�P���l{xfo�MDo�]{�?���W�c""�#��v�E��b3�սUZ�}�����ոT�e���J4#��72pEMc�zY��n8�B�i��r��"��>{�S�>��������ˆ��#&��V�E����|n�'_��x��,�s�޶�Ho�"��������n��xTͨ��n��Â D6h�Rʁ6���2p�|Q�$q�I��o�S.�
x�3�bZP9�t��h#{H)�c�,LV�i�G��0h)V��[څ����a���wʵK_�r=M��/���_WJ�D|��@D7�_�t���?��P����S0�#p��������`A�aj�Y�Q!���T'4����&�-�&���L\�x�txa�PدoPl���fpp/\6�}��Cg��r%����lKVkk��P�C(�U3�����1�� ��f���z��P[�N�1��e|���N!t�d����Mj6����@�n������cl�r^j��3�6�)S0�u�>���24�͍�[A2W