XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w��'���Om�>fp��(dN�?���(Tń!�+�Q�+��S���zm��Tǀ��e�Q�����0���=
ji�V,�Mn�$3Gs��l
��
�( ��=�	�~;և��aK��+L�_��g�<�y1�x¾�\�d���N;����i09�4�<ǆ�$�)����>HC0�Od2ͅ��_����)���0���v&)i:y�`�uK}�?y��35
Gڹ���u:�ն�Ro�r5=�CQ��qP��Zg��g���]�!ŧ�	�k�����s-:���F&�,����:h$'�J~iz�I��Ɯ&F,��D��R����"
�6`�����;A
��$k�2c���B���9�KjK�Btk=���,S5�]��#�I�Ҧ�ޱ�.c�!�Eѥe?��VBW^X�H�I�����[�F&]�^������T�ZO���ɯ�I1���.�;Z�P��tv�n��%#̈́m;��p��Zf]4��s,ō̙�mǮ�υ�>s5�0eA���b��/��\f���lT(�ؼ���uk�3ΊKX��Û<���MT�tF�QU���]��˥A��%��(��h+'���)�`�U�_ކ��&��_�?	t%.��������lO� �Z��KT�5���D��ϥܑ���֒G��?<SC���B}g��5���=��ñH��ve��[�X�H"Z���3�ZtH�6�@��j*QN�}�{��.��,_t�Ɇ��h�[L	WuZ��\
1��F3����_����XlxVHYEB    41a2     c20���:�lem��#d;p�{���bq\qr}C�,�R�dH�gP����޷���#�]������~��t��� -/1��7�'u�Ŭ��!O9HЀ埙0~�G����I(_�:�?��9�0�%�ԋ�<Ѷ8����ɞ��1^bI��-5	-8ۡ7WM�;B����AC�K>iV=n=��.P��xcn\�"�C�{1ji��l����9��8��C����3�`ć"�0���_�����{6���R����R��]��*,�R������~�uH�hZD;�c�Z����~�/&j��`�,`k�WN��(�p���N]�V��?�X�*n�Ԣxj�.T�O�{e(��%U������9�9�B,d+&<Y|�I���e��^���:����$�W.���E��n�y:b��2h��f&�5Xg�ڂS���˻.�貵�� ��eF��=l�7�:t����j��Sm-Ю�iTf<�������A�+l��W���� T�`���va�	�9g�|1#=hO���@
��4©�˝S��\-��;e���&�J.��#�dS��J�S�{�e36�#����"C|�-���8G 8]��2ִa��g�2�q�Բ�n�I�&xA�Ҽ|��9iD��X[� x@��BЛ�?�w�����'��"�v8��;[V���A�{5$X�\n[?^��v�0��sQ���v����v�oG��~M��9l��ϲ��R�$z��y�pS����o��~�)>X��wf���f�Z�%��'=�)���f�5>�9S�!E��3�b,3ua��mt��Zy�_;�V)�X�c��Y�\�����d�+ݱܻ���G�B.8"�;��g#�>�صJR*����י��ϻ�tU�����/���C8�
y����y��^��аdh�T�[��⣀5^ڮ0�A�A�
�uݴ��71Hjz6o]K9�=��)��&����Y&+�^%��C������Z �)��U��Ɛ�Kc�0�A�Ϩ@����@��(�,ܪ++��}Kc媈]U�y�Ы�T�@F��eB�������_Y�-��9��#��iO�J��)Q�>b޶�ݰ{+\p��_���\!�@1�n�.&H�@�E��۠�*��y�����"<0�>%s���7�?��9���C��v��[����-=������Q�6��l�_c���0�f�&��{7cd�:>�|�t�质��^:U��U{�Iw���+%ێ�ֈ���TEh���Od�����������0����R��Y�R��q�������u�}V����>,T����ҹT"rd"��Pa �ve�sS{v�^A�֞�P+�+	���f�cF>�������ܦ�ǃ�=7@�h|�0�6g�FD�k)`�@�B�NVi�R	B��v�8o�9�7���A�c��/$i�-iL�幜 x]�]q��&��I�t�771CN�Ə9�Gö�'�	G���Uf����)���]���LѳC�M�x
	���R�?)uŲ7[��I�>],@�c�ĤXGN"�Yѹ�x
P�^O�֤��8�ȴ����c�;V/�1�x�jb�֭vQ�;��ޖii:�9�3��3��q�3+s�P�gͅ�珏Aɤu^ù���@ŋ�i����so:��Б;����r�tH0�g=!^"�FCjp�0��?h���P/A~�0�SʈST�j�z�s���ȐM%ݥ�����-u���"�T�?_ ��ﺏLh�lWn~!�l?&�FR��pe�b�9s`b//$�a{�x9���S�=�Hr�J�5WS��R�<(
c�Tq���8W"���:^w���s��|)ag��l��M���k�ȼjx��4��K#��e�Ɏ��i0�s��nU�Jߟ�<�#6��ɯ��?M\��=�*Z����|'..�f7���҉l��F피z��W3��w`��;A��2���(`ǁ���{��v{������AW���9U�
c���]5d4��@�{�.��� p؟ �{�k�S����� ��&+���2�z�Z.��6��Y��+��%yA�@˂t���&�ƫ�V�~����bJI���ai:���hOK���O�����V�K=UHg��ߥ�q�lM`@HZX�lmǠ�t8�f��R&�i�����$ާ�)�fnߑ&?��mi���Z���ѳ>��&K�l�Y�?���E��$�f�R ~�o��e��"�3�h�)�*T͝��RO	.��k�h9L�w�y���T��'��^0ډq�B�P��5�[Fl�Ԩ0aG����.�H�])�	�Ļ��@�@YE��j1��T&����������TІW"�[=�1���X���/���L�꨺�l�w�MZO;�z���<�aS�kv�g�ۍ�4N�,A�$W%�m�h�'�T�ha�ߖi�.���)Wò��͟;�Ҏ�$�?ۙ{��|:55%ϡ�o�%�E�]S��30j�I�s��� �]�7t~���[}	�I����{ �ꖝ�b���O��%���=]�<����-�����?��S�	��-(�D��`��w�Bp2�m͝
g�����LKF����up��l8/"��&�c�VSU��{d�2	(=ǈ����>�Eˋ��^\u(�D&�߃���W��s^�Q��R,'~�[��8��2��>o��c�|��R�ē���8S[���'�"���Iu�x�®м���x�9�t�E�;�n�����9HK{���#YDڶ�=�LZ�({���ƚ�8����_��A��ݥ?|��wF��ؖ�#���	���:�yb��06��1/tj�w*�j���w{qM�I�$�P��g��~����8Z4q�Õ(Q���ø\đ\=��݂qL���q��*�	�˓����
��xi�&���힙�=��C\��gN�;e��(�{���7 ��"��ځ�>��W�Я]��5V��Z�o�*�|�ln�����\�V��`��lR�h���L�dL�B/ݺ]��߶��%k��z�^',ӫYF+������ڍ���e_��a$�q�����Be���s9!�:�\�