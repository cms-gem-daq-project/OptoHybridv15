XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ւX��\��9$�ȟL䫋]-)}��z��j��>(%������7���.՛�|��H�#^]RٚY�>�H�HǊ+�`�(S>�6�1#�F��Suc�3��0��X�ȇ4�'��~p�J���y���n�*آͷ_����m�*��fzp�;\�HX�����B��l��$�U
gB���
�w�;��;�|M�h�~֊ڥ�"��p[�_��z�,�	!��!S�O%��M�ZW�(�4)��I�;�]Q���rDg^BZv_}�9	��Qv�&�D�f�,E|H����l����������]�����8�k5���[j�3���NYuZȓp�a�L�V��������2�)�����򷟷�p��#T������Kef�U{�f���pr��7��� ��^�ln?�A}W:x���{�m�_OE/��p�*�����xs���0Z�&T���Y6�pajp6����%V�
��h�1�4���#���zW�09�Do��}�c	��F���Y����
ӂrS�՝@ɼ�B�#�=�3�:b�>�L
���4�l��܈�Չ�u^���]�<[����S��d�-��aT9�2~�*G��YU��T�HT��&���`s3E,������3��$n�5h�����9��yИ�����J<�����6������ �<�ꇊ�����D�0�9ca��R��'*��1Xi��A|�T�����
�$���y�[��P�"���XlxVHYEB    2902     a40��h�����a��RC˦������M�,���N��g�d����{-���^x(�\��#r�*�
��@���LRڭO"R��r��Mq�٬u�WJ+`ɝu��bwe��>��_w�<(�)�V�ϫW��[Mn�Ҝ�}I�#Р�����oN�Z)�z��!�7�O��dhY��5� �@6}GJy��ȡk�x7�}+c�rshŲ�ہ� �;�S뤖&
2a����&�'����9�]���%N��9������d��AԹV��WF���n�π��Z){��:D?�@�Ϊs�d������!����$��&cƙV�Y�CB�<�HĻF��)��d���`��V���־�d���+��v?>uG�0n�:� Q�Lɡ��MR^t�t���ƌ(	Y1%�ѱL�@����Bi�]&��D�rf[���nd>/=H�b�[�Jσ�9*w�C}�w�)�A���=x�2L�����!ǈn��ҎF t�}�~�h�$ϰY��&���Ƨ��_�ڦ�TJfU�����SR����c+���L�Ȗ�{�����0��$��|L��sD��l+��f�Gs���Oqb��gP#GaB�f��f������g q̩`�N�L�~�G�d��9�L�p)�y5Po>��b�T��
�����=�¤�_�x�^���E�;@���0�ɩ4��{��[!=������~��y��1��n�R��T�i�R:���h���E�
F�v��ܢ�5��Ղ= Y��K�z�D�ԑ�'�vajI�������j�=�BH&9+�$�?R��k�3�� 5�U撑�F8���z��H؉>T�_߭moC.I,��������j��\�u�E�_6<i6�������u�l5nu1���D�T�-B8�7.��>YǏMC3���0�%+(=�d�H���3w	J�*�D OD�zx�0�j .���c����K?��j���g��,·�8���94prx�jicP0��{�j(�`�N��)��*��ƻ1�N)�Κ��ʰ����	w��<`�����C���b/Ϸ��$O�*�"|$E�0I�<Փ������npw�>@K$�G-�q Zɥ/�n�C�8�=���VW���E�dR� (��Si��c0�#%q�u�X��֋vIN��+'43�H�B`�g`Z2��p���s(�������/�8v)�5�.���2g4D^�L ��1�F���M��-��R�.�W}3nU���=A+I�&`9��z�;��� ����8�0T̣�s��1��.���YB��[!���8Z�0+5"S9+�M$��Pr-�O\%f�T��G3}�u�U0�6��f�Z��ȣ�:~9xq0�j�7/�SjD�U(I��@�(XM֘��\�D��w���nH�cf����a���*NB�����Tc"A�Q����[�� &�UxM��s���\�Qgi���*g�>ya[�����|����+�k�Փ^��p1ί8�[')h�g�/5�NV�C��ltEq;�i8zyq�R��1���\pp�F�4��y(�SVɛʥw>yI�͹k�V��]����욮�VX�JƉd�l�X��~G���T�3�O$Ҷj�D�$Ѣm�P�4�6���ˣ/8�F�E����a^/�_���J=5to)���%_JO�" �V"4� �Yr'�K�S�:P��b�����i�O��AY�"���{���>�; ݺ3��[3��W9�����|e@i�0A��n�7�Y�W���Ӭ>���r�����&�4��c�(A��#������
xxX��D6Ob~HFz�������Z܊nԯ���M7��YF �@q跢��	 ��|�̀W�	�L�KGެ���kt0ri�Y��n�b
3#m(G�Vfl����`ːz-��ɢ#����ʏvz�9��1wqܫ�س��fa;��.	'�ƈ6�?Q'8���|r&�d��:��If�{G��+?�fGUꗊ��xe�XE`G�\l�|��F��T�i�,�I(�7�~���(� ����țMB57��c~�J�\�4<9��d�N��:R8��<9��|�}�)�k�c�8b���R"m��YէQ �vC�ybnJ�c��v���m�%@H#��b�����d����������E�Җ�W���=*>GD�Z��)u��`3}�W5"��a0�V"d�,W��Om�
�x(��Ge���rN���wN�xZN��u7�3��c ���m�L?������m/K�M�����^h�bH/KB-ް���>�1M���@���s[�����<)���q��)FY�=�&��t��ٳR������V?��EV���B�	6���`���<5_��l���l�7-��Ò��"PǬH���sV�U�����!�y��U��E��
��� �H�����ot,P����gpH
0�1�?�f�W߭ʯ�R���^����jR�X5��F�e]*���Lg��HY��)����Ԣ�F6�h�$���(�� ��% "��g�����-X��jCx����ԗ"Ks���^߰�F�~�N��C��+�K�;�T��5 �~R���	���G�nN| ��t��W�\p1s��m�R��X@�jZUY��s