XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z@O��v� ��J�Y�5�9���V�f�d/'�0�w�����z�o�D��m`()�{u3(���BY�&�H�v/�}������..A7Ȝ�)1 �O�,Bi4�����s�/�Hġ��G�n/zr��Ѡ���ʹPǒ�_���Q�lg���fxk��j�^�e���N�4V�G?�|�N�5iK��[X+�Z�����M����]�{%{p��(HR�#�b������9/Af�E�1�%y���Ԕ�Y<����Ő��]�q2*�=����3�߬Nv�N���6`S�L O�(*@yc �� �&��Xr�4��+7t�<T�)]h�ם��Ch(��t@1E�:3q`�Ny��?��~��u���-r� �(*�ا �qU���րj0��e��1C|��yI���D�����-����ġ-�����q~�wD��G�n�o�	���s��?��`�6���~�l���X�)3�(�H��+��]�5�D֍���CqK����y�e�Dl�۟l
���	��05%q?�ֲ{�=���굋�v�-#dڶ;ѳ��p�P���x��A}�G�ҥlGZ&�ת�뭕�mr �����e�`��٨	��k��2���x�v`3�V5~����nNk����ά��3��ESM�Lg`�/�� ���}c9��0����i���Bã�2��3�0�r�QOl̾������!�0Du�xo�������{�''�����!iǵ��	�K%�XlxVHYEB    156b     590��L���N&��n��iI"a��))�pJ�K�y��Z��j�u�jO�|�I���x�	�x+�zVf
��u�Fc������A�)s)b�u���:����.�]�m������~���0l��ig��D�����j�$;�ZzwE�p���!uY7X��~�냎��_��sng�b�}�њ!�.yu*2��������xF�����٠��݁���;=ON����è�U�F���<����;k���J"�rh����!��+�=��$,Hd��D§��+(�����`�"�E����Z,>ʴ%+��G�#/�����b�}'�?�哯{&OK��ι�aƌG�8ƟJ�<9�+>p�d�Ozb.�_Uq��4���q�Kz�]�i�D�/��t����[���0��Q���0��� E�h;�n��;p��γ}Ğ���2�w���nG-G��g��W��ӕ�|r���"��h�CZ	�Za_�'�SU�ٛ�ؘ�0����$��������μW,dѶ��D<�&�SE�+��6�-uq�������E�������*��pG4��1��.����$�ሄ�-k  ��f��֭�umr~S�4�w�|�bCg����H�<�^*M~	�z�mQ���Ӑ�\s��Cͼ��S�A�T�i�Z�3��� 3�H}�
O��xԀ~.X>�K�\;�N�оt��k����uS՗�8��Q��*1�8NrQ	*��f���N>eh�SZ�uϠ�tɚc2�&]����.rQ���mR�|��2�n��d �RI�oI�Tp�ȀL�X�/GCno�)b�[/���S�Y'"���t9����e�]�&���y�dOVⱴ4j27X�)��ν[���ԩ�s��o-��g~�V+����YG�W̅����$�#�ǐ	wX&�[ymT���[x�e��i� ��6�AF���>�![ŘJ�mRuNy�4^�ָ��MT-�$��]�ZvjT�_l�u�����c9P�V _ҁ��۫��T����v�=�4E��sDp%
��_d����vQ��m���2iI(\�X}b����d��*��<R�H�c�A�&��ɬ����7o{X�6(�/�cܲ��ll����a��N����ق��d�d�5'.��B��1|`���'����F���J�<�k~�PZ���@N�~n���j8�%U�È�y���q�#�@=-��v�����Ϭ���!K�q�i1�"u+ǌ�'u���{��b��>��s�|������Gp�߷�Z3�-�� ��W�!ԁ��~V�ס�i��y�X �?� �
�ev�e3���8A�����E���\hޚO�{[����8_�	�B;[%o'L��-���b����L6w^
�<J��Z�^�ܪ��"y