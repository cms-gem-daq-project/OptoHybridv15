XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������X���,�B�v���}	��{���Ա.6��,�A�.~=���B`�����*�:� �̞�2���)�q՗ƭ��<ѳ��յI����L����C\�f�'�.iptԖ�Xg)d�XÜHbW���	��L���	�>a4���t��E�$�����}�*�%��=�Y�'�����͍�~��њ�B�g�B��[TGC>��jU=��G�8��_g�]��T#�p��IR��%�	�T8�|>ʟ�<Me�@��(g�=��a���B�?�w����OP�?�[�V����ߙ����r�jJ�VO�&L$AV\&:♖�\3�S@�:��� ��̑�-�a"kQ�'.E����V�����A-��f�9B ah��W��g�BE���Nm��d���/nM~"�x}F�k>��:E(\Q�|��*p��(���~\��lvϬV�'�_�?6�'Ͼ������3�N��1�e�_��6e�O����������(�I�Bqu�GTh������(�t]��]����s����YE����I~�>�}sA�S]����YuQ���q-�V!B�[����8�D��Q{{�3��H^#F���=�8Q�8&7�ң��9�Dѧ=J�+AEIo�d c�CeP1�FH%��x
���E�K�+�bs�4H���{��/��7��ɔ��L�,X$�{��;�;�c��Ϟ 0o���c�n�K��{u��p�l-�ǈ%W��l!�C�H�e��oG:�D���)2XlxVHYEB     b05     370ZDaC�%C�TO)+����+㿽^�(HSńנfhzoZv�)�����#�S���t
�1e�� :$ՌG*�8�R���v-d���t;�*�s�6F"���J����8�.+��©�HࣝV����k�m�Ҩ�f�ʨTT)������uA. �=�һ.!D��^�-�ug;���˄���c�J%�J���ϰ��<�߾� ��\�?իV�s�
Qd���%SGc���_�ո4�9<ͧ$�p8��X�Z�gb��<N7��,9��܏X�7�a�`O��,�9�%5���]����.{�[��@���<��^@=
PMߧ,����y�3��~K��VugS~A&����q�μ��K����\k������p���o^�z��˱==F����(����j!Fw-��VB�w�~�5��;k/('o�k~g���A���S������թ����c��*c@�׳��K:D���2��˫��� @[��1W�a�ʎH�
ƺnǅE�q�χ�j�,��z�k��?A�C�|�������ls�[�?T�'�a& �>����B���m?���u~��v�+)=�ye"o~0ڮ��ԗ21i�s.����"����U�T`�D}C�.
���e$�n�9��z��M�Fo��h�B�8o�p=3�p䦐����G�E:��_s�M�h�>�.��{�A�m{���xx��S��ܤg���vf�O�P��lcp��t���F��rko@t��G��n�����ѳb���g�A|Y��/"�U�B�lMd5,"p���(�@M���`K׻v�=>�
�q��o������|ڐ� �>�[P�C�`8#�f^�g�<