XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k�J�,��M6l'��Q�F�������LmN2eJ��=Z�y� W�o��n�1S��\�����9/�W�!az���m���.��*��;H��zmJ�����p~o�E#�S<��]�#�M�Y��Z&EB��+�Uٶn���azj�kU(P�o�y���Uū�J@әS[PM-��\�����EA`z4�ݮ=��TkȆ>1�T,w�����&����ݤ3�Iu�%�?m ~�gY����1&QfL�oa��d�>���>�� ���$˻�%�$*{�t�డ� �I�m))���[����q}�G~�&l���7ߝ��c)�q~h�t��MB?��Uj�0��B+D��}���C�/���3�Dm�ǧ�D3M6�����CbKx��Ԛ��xM��"������(�w�UZ�(���i�v�7 a~�)F��0�a�,: ZM��g^"!7W�ĵ�xO"<�W��Z���t	Z6����Cp�݆�i�Ⱦ���̹��Zqܧw�.��|�K��b��|��o[�ζ�������pn�'ܫkq�>՝!^�ʉQ���ֻn��F�#��z�	�6q�ۃؙxc�������qʎ���)uϑ XTr����KEĤz�6��9�Oa��5׭��r��1�{��n�L=�uX�CnB��{oI�RC�&��1��
3� ��������V+T0� 2_6���"ӭG������ �
rΫ��zUB˶�f�iC.���ofi��N��n�DZm���X ϖ��rXlxVHYEB    1cf6     790 :x��%{,����h��V�q6UC��L	�V	E$������;e�%�I5�2�I���[b ���NU� �Rw�$ ��<��8���w8�!�����R��bWLs����4��9:Q0�P�O]"�m�N+D�)ahA�
&YU�8��s����z��	)�U�QF��*L<XB��{7��b
6��O�E@M_�s���n�m�ͧ:g�I�yp+�,������gl��5�y�B�q ��D�@g.��z����,�\��oro!���c��Y|��o�3bO��Y�_vl%s�wJ�~+�ސVP\�0l	���� ��<3~�I��n.]���]6�
r'����8�\ǉ飍A1�u�J[������P��M��*~@K'u�t� l�Yd�M�>���I��T�'��u� >��DC
~#W�&�����gwj���r!����^D�Z�}�D�	�/�*G���*t� D���)՘�}��)d�0���-����Q �ܼ,�=��nS�C��3Tx���L1��i�ރ�-d�ą���>Ȇʿ�߫���&_��+t�֚�থ�;��^J�X�~Ԩ�El��W|��l/p�Hf*��EW<X�OV��;��%�i���>����IeO�>V����A 3��1�S\S��>	��z�8�b�������~����6HlB�=��p�M�n�F����e��M��.��/]�ʼ�%T��ɋ٠�(z���j�X�!�$mF�>�d�l(c8V�4��𜇦"����[��^	\��k�۲����;��Z�l�Mn!e�5�����J����l�,���pu._���l=(�'N�M��Ue,@⣫����9�a��'�6-���(�f���)ߤ)����s<A�gXD�jpԐF���W���A6�L��\������穗s��4}b�	�_���S�[%��"�o�i�G��2���0��/�i�1ځ�2&�J~c�`y��T��v��>��"s���!�>���l�s]�|�A_SN�V=.+�,�Mg��YI ���&E����֫��'x�x��7��^T��&[eV'3�x��	Q}��>s�#��M���O����y�.��~?ڑ!����+W�Jw�l��ǭ� w� ���Y���^��s�̵�AI�f�V��=�IP��9.G�?�f��G��d�L2�!�+�.�p�!��x��M�7}/(d�3w���f�.%PF��GaB�b/��_��ǌ���N�p���x e��K�o������d�#�cvq�����1��j[�m��2e��K�M��U&����V�fb�����P�3S-�d����B�dl9�O`%jm.�#���K7q�,���L�g��sQXGrS��$�֯��CC]OWڟh���|������;@�(\E`��_�
�t��.��FD��'s���d<�sI���I�:���b�?ؾ��$����ŭ�u��òT�r(0�N��P����3ߒG���s��(<��Uo�QIk�5���h4'u&l�#��d͗F�:��e5w 5����D:�=��SN'~AE�HM��A��h����i�OU�^����D�8���J�oK�,I%�UM�t��L�\��!�V�ܻ����<��b}��-9��AqÝ�g9� +'�����*�i�ݴ!����'k�E��~%� xű�7�"U���u%]�7�|q�S���?�R}�}V�-I-��Qg�iMRi\���	�1��|��B��"�v�t���8���'�BJ�O
3UKU��#(�]�J��K�5�Q��cZ?ѫ�Jݸc��<d_��dG5M������h��g���&�5��m��|��x���ҥ�M��E="�|���!��T8/؀S:��ٺ�*�yqUxvt8P��<R���7��,~�1��