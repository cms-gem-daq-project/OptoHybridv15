XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���^�%�ء��c�,jд��Qc�����EPW`w��g0����K�3Iҳ\5�=���הNi.d����D��(.5a�r�c�֥a���U��u���_K�rԠ/����S\�K6w*,H�Y�lWq����v���o���9�-GƏW�|^Ų�!?�D��"<tȼ�� ��_1U�u�*�f��Ǫǋ#>y�q5�����*mIWP$8y�E��7� ��ypIgn&.lݷ.�3�[��o��u������A������^,���nR���y<�硫[�-[�OG9��v���6�2,}���pns�NG��5)����æ���!��m���hڪ����$s�1�M�-5Rj��N`1��HGA	���M}�")D��߶�c#���?&:y��ջ(�^�|i�S_#ZW�"�]�?Ɛ�Y���4x�\jono:Im�<�s������u&�|-/���A*��S� &g��%Y����n����c؎Ʀݵ�f���y՟�Z���&Y�ò?�@�S����v��q�<Q�����L�_��((�������
8Q�E]t6���xl�0��jd��?�=���|�5�����f���?�vȍ��D�k�P�W���<�دf0m5�����G�*����D��ԧW��u��U�N�(��������n毛��߸p��6��X\�l���Q��ы}�Y����#:����W{�Ib�]�#�S,�Z!؈���,^gZ�XlxVHYEB    9944     fd0sciSV���S�r�&|_�p��";�U*����9tEz�>�t�ÃQl5܎-%9��|w�����7��F�Uh��G 6g����[��Q�<R�H����굘�O��L�O،�ilx����U:!�B<4#@ 뤣�+�S~���Q�����xo������=Z ���+���3�]�2�r���@��"�"3�\�~��;25S�<��Hϩcq�Y��^2� ?��w)%?���-�	Jq.�T�or�`
�V��6��/6�r�ڀ�%2,
�1����|�/��Y��_�F��pEH�T��?�X󪩹�,�����3�{崄n����B1�;�:Y�g��0��-�\ULBU����ʗ���$��dm�� �<0�evX��tƄ��p���<�`vG�Ԡx":�V7$ǐ�($����C�æ�m	��)�����G��˦�~�iQ/|<���y�"p $G�޼IX;�|�I��'֝Eg䃐�9k��P�d+-�e�A? k���a�$h�XĜt��ܰ��~֐�"��pk#gϷ˰��֢wd\�m�(�%}����☆8�`j|�:�Q���z��QU�=f刵93K�����R Y�%��D\ާ�j�,O�)�S�
o�*�d�&�$N�"�mՓ����'f0�#�3�(��ZS袰�)� ����h!ܩ���?j�q}�	�l��W3�����/�`"yAM�B����ӵ
��})����i?��Ԉ��蝒-�XP\�xЦf�����:lւ�0�_<�)6���LfS�x_l��p��\�:��i,UL���g����i>��,�D�{�q. ���3^Y�����9U^J�f �:�,B��SL[mY<" ��8�O�� ��	J�|�Ĕ!�,�;���M��R���@�Y>�����a�밋���$˱�4�Fl`�����ʼW��݄�R[j��O��gWɮ�w}�EX�w�i�և�N�paE�#ű���(ǿ�|�x�!�{�
���ߋ��w��`Y�ʹ H��KG����&��bV:p88�d��������J�rr�8)�/&�
� |��M?$n�1{������tA.���sϚ*:�d���Ś�%lQ}�[3,�m�ė��ɸM�:�N�&�̞r����RX���*ɷ���'#>�_�
�� ��EarW�̓�:��$L7pQ�Q/P2�5cM�*���e<���|> �X��n~�E��TN���
`"�X��4�P�A�Z�\�,����7���dp��{�o`�!<Y���Hd�ńۅx���_����H޵A�dK�����5~◷�����x��ײ�E�6�ʴ�X�q�+J�2�L�(#SY��� �����Q(D��C*	�)T�]�a�
6��"�-�/[�B�q@*��|Ѱ�v����9QQ@�ix+�'��k��&T\J,oV;0%4{O�	vwE�t.����҈�z��|�n!	��8iE��[�[ߜ�E�	M!��6�=�ACUp��Tz=F��<9������+�[Go!��1�%�33��՘:~*�4��ļJ�-�ϊ�F����������P�I��>����Κ���q@^�G�~��c֭o��pB)������K/���/pqV��;O����N�q0��eY��c��n�w^n�� �8b�����w���[h>���j�;2��f�z���8%a6O'���s�>=�[bT��dGt�A8�@ORg��y��AS�������3`D����t��a��,�BGO����p��g$��Ep��]K�y_�c��Wy�X��FI�H�(�DnA�O}-t��ڦ��C] 6�*��8ُ1*H�BA�1�]��e�ˡg�2��Q!��$��2�%���yp�Ԃ0�`�ۛ�DgJ^^ ȔSG{��e0���P��_}I'�
�H�S��xts����m�v��]$��1tu��YG�%�*l�y>q��*$Шp$\f�fF��U�����'j���]�}G��������e7(��#'϶.�� �Dt
�� �9~��0c����s�Z��ͅ��w�
�������T�>�VyK	��K�F�5
�b�%�`�r��:��ߤhp�h.X����E�A�Fɟ�.��Gi�<��\*^�=C:�P.��41����R�H3XJ@�o�"���e9�=��|�X�tِ�Z;��u9AƋ����ԕ?������1��r��G1�b�O^̻b��G�hTݭi1������N*��ˈH��z�}���w\	�q��	�����T�*�s��]�7��p�( &dr'��&�[��0�<��j<jM�Lě'�����G����eˀ	>�Q���LF�(�[� ����Jl
ٞ�#\P P孽�I躆��Nӂ��shy�u�v���E�Jr��/�XX����y<j�˦h��+9��qz��{��B ��F=uQ�E���p�����-ߎk#�No���(-����SC^�ؼ�n���Y���� <�A�����Q��0�F�uD�aq8o�����t ����V{|y*V^
�~��Spk�u��u�nt1	���K9ѩ��4f� �V>J�M�����)�C�	h�|�Z�c}!��a�(�����{�H>õ��R^g��tN�|h��!�:����������� �Q ��]���GfϺ O����Q:�_M+ҡ�.DB�9��W=щW��`O �D�]��ڪH����:�+���緡��PGϊ�!(���P���\�D�M����*��s�i��3��2��(M���5@�6Z,f&��;�7��DmO�H���1�k?����2N���$P޽�ȓ�@+C5�
�|�4C�i�iB���4Z�������3 �@��|űn��}Ijӱ&�.@�󛅭J�5�#\Z��#Ϡ̐������+D@�}�W0w	���g�~A��)!!5:���1�dgZ��T]X�v���������o{9X^6��p�ܬ5jj57���K�fK"��D"�Fok,�O� ��k=�DN�Xk�fn���k�
%�Ja�I���Ө%R�[�r{�䅣� F�����t��P8�͟��*�sa?�
��xX�gZ�J�����:�&a���c��Z=T�vE��{In#K����E�̀I�<P�S?
I��� ����չ*�Ov��Q/n�ј�V���V�P�+�Nq"+��%�>[�b�\��7�ї�@�.�B
��Tɏ�ݪXF��X��0FhU���:���!�ω����Pө7�82sׁ����r���W�n�(�������"�gLgv�^֮#�$���F+�_fW!�Kv�G{����>�}�?'�a�oo\@{
b'���.�*��ۖ�����%�����#O���L�:8�u�(q?��|aJ
��fʟ���0ln~��dM������>�_]Pf�bA��CK�s-�bsڟ�GB�[&���	N|x��ڲp��9ق_�f<�<�����l�Պ�q��"Fc���G����{�$�z0Km�q��#X3��dAl�ǖl����ߪ����~p��VJ�
�mי�o-�)U�C���b`�������:L������WW�
S|�^/>�
+ӌD��8�.����=Z��4~fT��M�a��$.����Yb5�y*���<�e�.�?�	
�y�Y��o3CV�Z�}!����{����zCp�n~`.��RU�)�]F0)%+�����U-I�(T«m/(�)�gd�Sjl*�Pf_1�`"��+�v`��^����IE-�<��b�@1J%~�}4N�9*qCW�e�1�)%�N:����jq��E;;�l#��|2��r�%̽�e�UI1�X_M�3&LW���۱?����x�ؕ�gA:Vo���m�xv���cx���_�DT���($�]�Yd� �j��j� 5~�����=S�ˁ���"۷�(G���i��	�K���B^�q�����3%ĀTծ��02D8\th7