XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�ڲGLޙ۸��&��p��i'��s�N�s��,�3��+�I����-�d�X��Ls}���"�_��O�6�CUvl���0�s�V\�7�1-�zIHi�\p��9%<��?���y�N>9�ƽ��'�s9q�8�!Ek
��Q*�/C�V�����$w%��(^�US�{磒�C��$�WI�Q!���!p���	�'^J���"�QQ����9�h�G�o�5�zQ��y����cVb|۵M=��hJ�o{�@�8�0�ՑCU���q��N~q8�WDS��3�b�zpYP �_m6����R���n�J,�O�c��D�i��G��V7N��	J��t�u@bm�ΰ�I�9$8%���@�'��� ���/ǜe�DQ�#4e��P챰l��1s5�$p�Y�wpPs�?�.?��A���1)���P��kv+Q�gI >��<����l�R�ڮm��p���O�:�:Go�-2�n��,�R���wLV�)�h@	��p�lBJ:�
�܈��P�V.n�4C��� k�3S�K4��w�`!4,��}b�e<N����6��&?�� ��%��Q�%��RWi���D���O"��;	]�D`�?h�����o��{�xe2ǟ��k.�J���>��5�%ы�2�$���<���X��ܚ���?�ʝ�c,��I	��Y<�ߤ���+�JYħ��	II�}sطB��[���?e�=��Q�[���j0h5��TJ��_c���XlxVHYEB    1cf8     790A0���W% { a�`wV"2�S^+xr���P%��|"��H} G/\������ZVrI3?�����ٴ�f�h-�X���M�F�Qi��CPr��'����P�����`�O�c�Hf!ٝ�{�٘.��v=��txp)���U�-�Z�i���P���J��Wd�5ո�c����6�#au�pA���v5����ҳ�&n`��7Aۂ0�ӿ��)DVY>���ro��hY����B0��N"lS�%��N$gVr�c��b�ئ�;�ӆǮ�πSs-p�?�@~�eL$�Bh:!���'��.W�|$�폤��nH�<w��p�5ޠ����2Za{e'f�����ih�l2��o�S��ʲ֧M��j��	��n h��6;c�s} ��*��X=Кw�8v�xqu�����Z0�-��>DZ�!����g�&E�|2QdZ[��yk�T��j�@*��-�7�!*�Y����;�w�0������ʫ�'�N�i!Xl��̘�˧e��.�[�����K7�ev\VA�L��N;�����n�������qp�q0�6��l`I��/��ߞ�F*9��CZ�M�%����eo�L�\��  6ڎY~?N�4���2;���g,ma�V�4��O}��2�����dv�# ̅�1V���_!h����`,\��Vꨞ�-��|��I\�(`���9[�������h���K��ݨ�= �s�C>\W���4�pؿ��K*
���4j���6�:z� �w����[��
o�`w]:d��V����(��|XZ��m���l�AI,���P;+=I��Ғ�Q�OR��_�Z>�bMɉ��M�G��ρ�Y�����GG�L�2��X�?+�?	��{b_/&-Ljo��!�!@����^�P�8��h���CI� ��/��ʔ�v?��#����g�����ey�Buna ݊����=���'���x�w���Q��kfc:���c�9
��������A��gv��5�1��^Qd���V�U#�5�x�V+͕څ��v8P�~�`�5H��\`F\h�	�*�a�\����Ua�L�DF�W4[�C*��{{�F�u�-�)؆W�<K�B]�tO@��o��B�i���۶2�_I˕��4�,k�d���c�3O ���0���YÅUrHn����B�f����`i�JLjց���.x���T;��'�C�Q��^/�����:չk� 6,�wޓF�%y�������yIǂ�Ǯ��^����LQ��B��re ���D���H�u�K���� �9�3y�-�,��|��H��ũۂ�w��:6�Ʀ����rxv]�d���fz����:ln6�	��g��Y����^���.��ƿ���A"��F�҉A̖�����Z�����	���t��f��-�#�9 lW�-;i�'�|ě��M�Iqq*��g�u`�-�]�qy�x���홍���j ����{T�GL��'x�Ѕ���P�)CTo;���`�ź׃�������Y���i�2J�m�-�j�(��*W��=���U|�`����H��D?R�����G.��Q(�G�5�E!Λ:DiQ��{�'���Q��b�(�pWG�K��mZ���G9��l�	i_�>G̬��řd�\{�b�Z��l�x�$��R�9��/#>�H�87�a��?�!$=UoH���}�.V�l9)'�Ɔ�%
��#U|��Abp��\�P���]�i� ֒]���uF>G~E������p����H6���Ň>����d䁣rVuY�Bb���t�*ϋNzT�1n�'���1�nBhR���m�>ޡC�-�)ti�ғci�IX��]��m%���/��v&Y_|<M	sN��[Vݏ�:ٖQ�,�{GOC