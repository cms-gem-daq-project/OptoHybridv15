XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����gg�+�ړ�m�Jk�^�}1;������>�Ķ\�U�&��M�v/��_t�c~�հ�D*_'�A���o2���6h��c���ݺ}-���9m�ډ�<4nRC�J��r���B&�������~&G�D����}E��=!�ĽX�m�u�?@0��q�3�{��kU� ��(�����}�s�5N3*�ҩ��6�cv���Z�ȠR�[@�F��c��QL���p	��#PN�fC�[k��[�J��}m(|u+w���w�
������Y�Z%
kK�T��ema?!`�vM�~�A�U*�7���]�>���|��8��w���1�[��?n��7t�����;�i���/o�5t�: )�� ]�
(}N���xT�2�7�@��NI�����8Cv��/�l��HYB��J�ϑ��N�.q���0��" M�Bč2��"��
}$�ܲ��_F=�8A_j��$w�����oj���V)IA�%D�0��K%�;�yhKG�	������A�_[6r龰��M�a�N�Oec���u��j�07x�ed��v�����7���T}�V��5��0��cx��{��
�JN�t���(��MN�~�tY���]�[ɴ���n���fqwdO��T��2���蟋���Ql1���f����7������M�3�'J�x�R��y�*���Wq�X��0�@hx����~���F�!~�i�G��>�Ѻ=�m<�HR����4;����7c�`�庁R��5*���XlxVHYEB    225f     610���H�V+�Au���Eˏ+��!��ivg�����*��<���lI-�lh��Zz��Vͯ�RS�b��]����/�$��� Im�ޣ��]�_z*|�t듛���v7���Ι
k|:fR��M�P<W1�� ��,|�j�W��.��_J�d�ި��6��h�J�Vy������1z�AE��Ĩj�1!T�n�RC�)���d]w�t�#Xm�ɝ�ȬR��:�%SX��l�h$E�j��m��](9�g���#1;��)T����F�`��5�w�y�ń^[i�D`�����݆�vShOǤ�j����9=s������Íi�˽8#����n\�:`��I�\&u�xR4��s؍���6�e��|�⾞��N���_�ՠ�k��U���5T�@����:�|�h� �ww;�*�j��

���<������k�XZ�ݒU���]�+^� vEw�R/�ѭ��Ŭ��5{<Q��l�[��J�����T�7s���<t"
�q�>�n�f�S�H�֏�7�*7�cE���	�Ma\��i�c)�J`�2#5�*x&j�O�YwI�%CR`���qa�'�}����;e?��f�W  �KYѧ�J"cB\���7���m��F]�I�W�����<�n�Z�@d1q\8���f��+�Z��\���V�춄�&��</n�B%��#�sc��]�.^��3V���*��`�`&��~��q�J�_��/ r�Hߚ�+���zT�j���.�����p)���E���2��o�����[��lD/��p���hc��8'륓���ӟ��,�<���%�`�{�*��b�f�4s�B҄��5a�o���0��0�n�����2il�Rx���֩����^�	�3���j���]^���Z��6�"�H�hl$��5'�����A��S�w?\�)�����n��Ek_0��O���������yHKC�Qv-D�)u>��h����=��
�""W'�\�qR�����S��+�Z<K2�^�[qۄ凚�@�D�|������H�K���WcH��o��\��E#������w�I�E�j��/���jA�N�[5|t�O������X��>��0͹�RE��Ƽ��'�ک�/Y�,7�(��I��hhZS��p�|�N;��\�jE����\��M��Y�$�B>��� `��0B����ɫT�5�{8i%�,�X��B-=�f8�Ums���v�KBg�QV�1d���TG(����zFJ� ��b|�X+z�~US��Ҷ2�����F�����n�o5b�M6�y��W�P���1n��'���~�PIy���^���H-\\��tV����:��������/=��Ɔ�W�N k�V#�T�mKa2ڄ��t���L������U�A���}q �I�Gb�U ��ĩ�r�=�~Y�魞���)�L�7���i���k�h}j3��_���۽��q���-����r��
h��]�v*7����d�)�F�1�<xS$�ʏV�V2����