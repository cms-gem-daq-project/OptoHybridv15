XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���r^��֖$�&�I��6\�|�U���
��yWt����=O��Б4��F��1SV~c<K��ߧ��5k�5��2ȳ�7@_LW���,����L�:Q*ؤ��&x%l�jq:�h���s��$nA��"\�1�V$�A �ɒ9��{�ib��:π�sd>�ؠP���&���*3~7#}�({4�I�~Iąoq~]���@�Q%�+�>`����Rj�yW%#��E{��z6KyXߦ��<8ʏEf��1� ������6��9eH�X�Yt��$O�bv�\a�ӆ5�E��,>o�>|C�v_9�P1o�ZzjxǛA%F�mk�
E>e3tK�ߴ�vr�9�F���k/ğu���*K�YIx���ݡ��.��8�,�ŇX���mᰚqÉ��-���]���w*}��w	9?!%T�U�����Ǎ7㼛�8��c�?O��/�����/՜j�e�� ӕ2��2'�)�|p�5���~S�R.,s����m8���P�(�g�eE���6�!pZߴ���Z��Ͱs�v���@��b�����\Nw������j-m��@�F��M̽��H���,O��X��r ����f�0)R�"��NY6?"��	L�Y&����)Q�z�E	<w#p�aN8��ć�:`'<�{�cYn����,�A.����{��	��HH�|�s$�x����v����LŴ�۫��g!��S\��3�]����<�}���ǯ���.Sf9��]f�,g�kXlxVHYEB    5ff4    1040�I�u�;�.r�����d�οa������|�쮅;�l�s���O����U���\� e��g6�1/1&��"t��^sT<yT�A�K*|�W�e\�\�	B�"����&���{��Xe;L4����W�4;P(#vr�F�����Ӊ��z_�G�E+bB�ׯA��4
w�'H�9�{���`�|�_*y��M~d�ݚ"�^p҅gfR��T1|51�I�$��6?T���_�|u����XTg�T�c�m�i�qțX:�3�_L)���Wr�%>]G�Y}�2���ڥ�.Y�F���v���Z�n_`3�1��:H_ �!�u��<�@˃��c����fLCKѽMb�|a���+���{������qŲ?��l@��T��M��Нb��pv�>с������ƻ�S� � �	^���ݣ<���e�����ti�2'z��>�Ή1�"���7�c�`ޅ`�B��B�ɋ�S�z�]q(�I'�6�E�܍Ĝ�V����:F�~�L.����Θ\+h�4�9�!� ����1���� ���?��P:���+p�ɡ�~��8�I۠h���#�?���}�%�����C�5�I�P��*��G��J�#� ��ds�%�c!��l�T���<H��H㆝F�j��!�)��I�9���@��[��;�t�^��<t�:��;���	UCU��`�ř��q;L�,�K��V���Z}ƴ�n͓U�?��5�h,i�~�w���[���)������?@7��t��;-��M�
���y� 4��Ccb�K���O�)Z��Â��&�Ч�R�=~�G�e��� �U5���+�4�.A�ϳhY��)�=��|�U���
ەHgk|�[��*��6������ծ��cP����i9qW
��ז嵐<T�u�c� #��$`�.Ƽ-��)uզHߟ��>4�4�aB� p=��x2m

+�֕�R0)��:�)����Z��	.���	C���!;#h>ޞփ-�3�s��}�`ꯀ�܉4}��Y�k$����������)�Nlk�uWo�D�Jl�ݗ�5�I�(z慃��|���v�!��&x$�(R��������d{#�4�e��cp�ܷ�Kv��؄�s����Y3��j^���"�5v�����Kc�����T%�A<U��W�p��&�nlmX�j(k>�N�m��E�l�Sb�luВ{�Q�s��Ӌ]|bo����Ks/6�{�T�U6�@~A�W�����d')Rch�9����>�S��� �_o�]7wV����6����cA��X
�cD�oy��_�x�1S��h�"ˏ\��b���X_�5Z�0<3�$�� ^�*�i^@�x�0g�M�]4'hXEY�:�Q�:Jzb~Z�r����w���M�7C��^s�=�8m_|.tb��V{+$!9��a��t�����@x�b��kO0�<)��]�a@�g@�Ay��	3\ӡ��~IkU�r�ӪS�x��l����e��8�sZ�(����,�.}�Rz���Y�B�Gz�^�#1_j�%�6�:������+�Dp��JK�0B.�2q��}����"y:��=�x�]W��n������U5nZ$r��ΎҼ���;�MZ�h�ӓ�������㮢�U(fȻKy[6����y������k�����1�x����C��qv���S��"˛h�1�J����r`��h���WC^ٚ�E<��6n����C����P��wo:���|�e���?.weH�\������~E�g#��>s��^���O�f�Q����p��{as�ʙi,)	\�cp{Q��o��=�qY�@"ka��0�Y�4HM�=+��m��1�(��Dm��ȼ����Q������'�"L���*�c~�L"�6y�'|VƲ�$/��^�
���A�t,�CZ���Wm�����x�I��I;��Y����o���hW+����2Q�!��:�2*�)}�
�Mj��m���5��CL7`j�N$V�ڀ��;(�9�{pB��$q2X�YVK'ʫ����n�*4�#q��R��b���o�c�\D��I ;z����y;[�-�a:�Td������Υ��? 9��j؊��?h��fՑ�Z���T�c�HX퍪 El����#�g����Z���4yrW�`��EXpr �7��d_�Ы�pk���a���/�8&���]�R�a�la�赠��Lo�\#*!˕���֕/U&{
�GF��ev�{�	�Q�`�0�O���6���.�Sx*h�,�f��E r����̋�q���A�li�-��A��Q!p1M�@�Ú���KC����
�1	���8�V�m7�R��j�����շg���^�B�F�!���e,��A�/�wQe34%�頴����(��u~V�/����_e��n�%P �]���W���˾4SB���_���2�?��4ӣ��iS���F��8�&_�a�ۛ���x�w������=���k�Y��&S[��NK�Q=��0�7�03��������Ju,L���"oOj��u�|�7}��O����⯋��y����=D�0C��<��v���)�����h9B����U�}�F���$�	���f�A ~���o;�owϳ���]�����D��I���x��C�1e�E�;OF�f�����ą��9&v�`2.�=��ƙ�4:��؍�9X�4U��
^p	���Lx� ���s�`����Ga�>�����<)���w�/�S�X�9A��'-JZi}W+�tX^��%�ѝ�că@m+���v�2QP��g(��7���##u��m�^�T|I�L
8�S2�Wtp�F���=S5�U�~���D��������
��=�;ۥO�a�E�Иg:���"P<��49�R5��jE�pR�����W"rd���m��%�˰�Zx�XH@複dms����/h�E���P֮
��q���ɪ��D�@�B��'��,I?�$}dh�0�l�Ej��m����4�k��}J��t��W����#a#��Q��,S���Fa?�))��=����<�;5���ld��(�����l��UbȮvU&�:[���Ź�Di�x�2d�`�j�(��A
����G�vh\���BKHUǮ�����tnA���Ey�-�,�������l�}�~~�H�4H����B=VDz���ʲ�'Ҳ�Qt���o�������%pfܧ���AӍHz]�褄ךj�w7C�`�����N�#�����(ք/}��؍W�*~��m>�
Q4	�bv�A��P�$�ZI�"V;�{;'���-/޸I�?[qz�J��J��cp�L� wۀ����W�1���e�]���qĈ�o�_Ô�٘�'���0�)��ꛔu���QGP��8�dn��j�y�Jȑ������q|z�����~���{��\��H%�o؅�;�c�%W~��k8��y���Z�ܿg�v���4]��*vf�x?�(̻��ڱ�Ϩd�r�bH���&ȶ��r�r�"_�o�J��ur!>aj��Pr�:ө��;#'kid
���54�Ҁc�b_���B�C�483:He|�gڧd�4����Wm�6K��w�����|�=p}r�"w�{�!���%�)��Uߞ{X)�� �lЯ*�����`#z+=޶�K]����������1���ȹ�X�lFQ e�kD�ҝ�����`2��4� �+�kY�����@����I�¨@X+�_� *Q��>�\ �pZǔ=�g��\����Y�ֽ�^W69��A%F	U$N��c�g�u�{�;�����~�O��j��<	";�~��ݮ�H.L6vm�������0G5O�h���r:���gza@F��E�+MC�B�sJ�<���SP`|�e�/���q�p��մ�0��o���cu�oO�/-6��%{�4�8��-�E=#�$��
)sF��)5J��E���Im�4�|�cއ���R�?׾&din
��mA��D���eN	Յ��G(�$��E��ܻ�������*v�T8�p9|K�Ì���W���j+