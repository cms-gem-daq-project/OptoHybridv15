XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��07:!,�.zC���b࣢G�xa��ͺ���b�pDЌ$j�����%f�;�A9���c�H���OOA���楨��W��S_r��Pc�G�Zj��)A�;=��mnL��A��#! [���|C��{��$��E#��R#.'c���wc�@��b ��~ZXk���l\�ΰ�?5�`a��t��P7�x$	IT�C$ny�s���#"'��yBKn��J�'��`��r:�X*ru���������i&���=�����D��|SybH�=ܺ�/^9�f�qAet�q�za-M�{wm�D�ͩP�_չ�������_�x ��!y��E��ϵ�Bt{E���B��a������p���<{H�N�'����J���.�6,d����2���I��0���E��"kR�.-0l��Zg��(.�1�f������Q�nf^)K�T��fާ�m�p���
�nP���RՁ��+~}�����ky�w�e��%�*�?
�Ю�j�0[�����l�T�>��uB���T�c�_�$BRb-�Eg�N�tI�DmQ��K��q�0�Щ��a*b�|Ƭ��ܒ���:��/|���ԛ���su"�O��q&x�����0:N�/��%[������k8�q{d�9���I[_�ݓŵ�a��M�lqJ�̉�At6n>r]��*��h�f�����$z�����SI�?e�벓�p;M6}���MG��W�uqw�����k�}�� !>(m[�1ˢH��U�_�XlxVHYEB    152e     580B���u~��W�G4�����,��§l/:��FM����X8Vo0�C��e_¾��O��m�.���KMX+>e�J�è�K0!+�Ye�d������l&m��C�"\Ų�=��105���kOk���q�V��VTA��4	�B��#22�������̉�� %~K6:����^��Z��WR�'+E�����i��2,�|I}���T�x�+�u��P��~��g�T'�ɟW2�����c�ZEB	m%��R��ϖڽDj�=��3'� �,^���+�TI��!��YU: N�����^��O��M?mRT��mjP)�!���O��K��*Q�>si]Z��k3'�Zv���`��)�	V\����8�\���GQ��JT��~���Rgq;N���.@pPP��ܩX�b֖Y!ድP]�/��|y(�u�F1}&��L�!���/6��Nh����*�)�c�� >��
��Dx�e%��Q���PGq,�,�rt���G�Z7�'����NLe5�SyXR��M����(��g�:� �q�r�03��J��;cn���TyJ��[�/&l�9��l	�rsD$'��i���O1��Act����o�|���m�xb�v�O�Q���NQ��
�}�2g*�z 3�}�����*�\��u���z4���p�U�7(��(C}jN�r�G�A��0/Ͻ���K�\�+�����\�[��4�"�����1�n��_�ފTk;
��`b8�8ʹ�%���p�/���ι��^�vr��ܢx��x�����h�L'L��]����c����wb3��9��!�����=��R��7T'l)��i�ԞCK�w��'��uԬ���,�]�����V���X��_՜ G��Lƒ������,.S��"�'���'0�>�f�O�9�Ʌۦ�mF}	�ʚ���M�>)^m�^�v2��m���n����	��-����腊��:տ��_��X�j���K�u�����&6.e�ݸAZ_��8[���F�R$N%E�m���O�w���Gp?��^̦6BIf����� �h՗?[�8�`�JPi8�b��4���d�#I�m(�i�kHgy/�?��i!=��n�'��cn�*,W �%���c�x�y����W��j{��ITT4�h��'�E��������E�����ӭ�@���_���~f3eN��v�&Ut�	��
[�9O&K����<�3�7��Ӫb�;F�n�hpoY�I��q s�"��\���8[-�h�O��=~���E�%�"N���.g&�����S���"�[��zx�$W�jfQ�ЮNl䒡�����xF��L3�٤0�qZ�b�6��]Ǩ���I��R���R�3P��
n����#'�2�Ms;[:bn<R��