XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q���/K���Z�P�#���VA�����z���x|���DτiJ}�	�Dޱ���T�K��Vw�~+�Y�Ӡ��o%H3!˙S�pw��������]'t+se�=��=薤�ra�;�$�7�Q9��ZP�vFS!�B�Ћ�C��3�<�R����.	����t��k��4*X���Wk�|�%7D��)t��ﭰ�wun�͸�z�jo{b��;��Rz��S����}H�[�l��Quc��>�R�����L2ZL���������s�M;j\�t%1�k�tz�΋�we:I?��1T[�R�ik|��F��X���~[Y��
Y��C��q][,�[������'(��<��cb�=��ۧr�g�q�7��RM ��A�n�������LO�c4�^2��}�F�X����oHٓ�G��C��U5���M�1B�����w���=!ȏ�t��@%pR>6�@Z���Oˁ�M��41��N���ƫ�́��x�Y�?�.Q2l��8&�Ҩ;�1i5"Y��o�� ֣��?*����W6Rg�I�J����X��N�jϴ����XF���C�"�����ʣ�{���`�D,�V �]V�|oo�d�����gC�C�x�6��L������,дl	Iɑ�e��Ы"WP��}C<

�a~�zK��#�EZxy��EoKY5�L��r��,P�P��dz7�&E�/V�10SL��Y��٣S�R�m������ˆ��=R}[N�19>�	&+p� XlxVHYEB    1c48     560�Z�Eϧ?e'N�� �֍��FEX-��Va�~�25x�2On��hqkژ�+��D����!�أ�k��}Ȅ%���G�d����e�˔�EA��t�xx~����%��Zm�9�rc���=r�ES����.��kh�v2&é�e�Ə�g6--gz��*G;����c��f*��a|(X�Qq�F��f���ύk�I!�C�K��6^O��þQ�˧;Z*�x1aU��'�M#T�vBr��Q�op��c��?�BY����ݷ�R��`~�L���}��L�A�3{���[G�Ҏ��9F���2��'�f���ؽ��� ��"����gz�?�٦�*$Z�U�|��$mW1��1ec�S �C�M7?�hb�V�������]����<��n��p��R�V�A�H��A��_%����⑗
�U�7����XG� c-1�X�Đ��v3���Fl#$�<��.8Y�ϻ���Ȍ�>z��v��~׎�G���9h=<Ͼ
d���l�"���-�	y���1��T���4b����	�u�]��]��$1wrG���˻��Ȟ�ַsC҈"Q�4��~r&��(Ag��ۚ��v�?TI^� ._�=aС�X����h,�:B��L��g׍E@Adi�!H�1���FGMt؟�m����iٯ�m��2��yM��l�}3������V���M�禨E�����#���YXf;{9�[���@��mK�[������b&C�NfN��[ 6P�wn�@�ozq		�+��!7L�x��@��M���أof�q9A����+�@xG%1i�T�)��j�qH�yB:ҭ��Fx.�K�F���-3^t���K�BV�Oe牬'�u���A�:�)UtӘp�q׌�k���㦒X��{
,�.E��:� <RC�~J���0�5|]��nv���^>b���)+�i^f���-NmN�oϊ�gI��q�&����j�;�����A��xA�QW��Y��Ȃ���~�L^�z��%��oܗy
��[V�F���r��#6��.s�vչ:H��]��C����A�ô0Tk�i�;>�I��Q��e�׻Tņ������ߴM���꯽P�і�r�@(���B~�R�}va5^�=TN՞��	���INz �胗|��Q�%ZOo�� -�E��|�����4GK�ç���K����D2��Ѯ����t����{4�Fګ���e��xt������ݏy��T����9qr�)�� ��\:`�v.�+z�i���� ��o{	�����f��S����E��*nF�"Pd�|X����.��`ϖ��X+�4j�D���JG�ҳiȰ�/�TfB��@9���b�MN�