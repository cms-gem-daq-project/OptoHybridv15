XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�=���sK#j���	�#0߯�12�¶(!j%��b��s���̙P��Zh�Y�������h��U[~��J
2�h5������I�w�ȑzӳ��/2�ٳ{~7lV\�l-�����k"s�2*]��23��5ԛ��u�����+u�)�u����W��9��� �����@p�z/�^���FC'� K���� �-ŗ�z��[�d�Y��=*	T�4��\��]W��p�(�pjL潧���]���4�E���ĵ0+�JxzLSz��1xA��}�����]�x?��!׭
Ә��/��V�;�}��ay�� ��V��h哭��zbX�|�*F�G��<'�X,OO$�?
i������_��Z�?I8�k7$��P#*N���T�E�ZH
�jq�	�=��%�1^YN��s������!g����� ��w�p��q)6�U%"�2�9���8(�����n�^R���o}���W�eP�>���(kY�43�eIqM[��P32���"��=⤦��̽{�Rl-�uyX��Vf��s�I\���e���U�0h�u��"�&�hZ�c��S>cw�׆>�̑�S���vе��ǹ� �/��Y�h�xP
���C��rS�ڦ~�����gް~0�{�2�&���o9ma!Y2tO���L�}T�����@�J�B���(�5�l� �rrF����ǻ����X�M+HR�;���<sɻw1+����Kd{Z?q.,%*�%M�5���w�D^�qB�XlxVHYEB    1001     490���;0 |����#����P���S?��S9����D�t����LE-Y�鼺ǹ��}�V�h�ִ�<54�����hJh��D��7�3]z��mͽ��q����"�}�3�[{�����S���SA�sL(;� �������W��tIY$�͒˟�M��vI�Ne01���R�����O�T� �x\Bm�B�S�i<X�u��ڻvd��Y�2s��u�����iX��9%T}�DLPrͯ*\VT�mٖJ��Mf�'yv#���&�6��%+[ەS��<��1D��
x?���*��������D�Rl���>֠y��r��:xES��eמp3b;��@M)�.����k�����WdӣfB���]�'���AO���T�B^D�Q�5!��2��WQ���XP�G���o�fK��[�[Sh~V�b{~�jݭ���Ș�����Y�:f��mͦ6͐�9�c���6�X��Ƃ%�m�+e�s�H�ff#�%F;:�8����2H��y/���G��L0(����9Tb�kgm��}�8>���Ʊ�Q��s�� �drM�n9�����~�K�mr�'�e���c�L~A�C�:R�.�>�??�x�Y(2���P��/+�"Zj���}�a`���b ���v$��~�������We�j��}�y`~b��+_n�
�Ӡ�Z��hLb���c�y���o
9��3/?�@��:Ϡg���I5Urx7�PT�ҝR�T��H�A�~ ��e�k֒�2�T+ji	^��S����o�;�@���]j�� ȦN|o��d�N(w(�п�M�{&|K���0~P���3"�%A��qk�^�w7�����A���o�՞�`Oobsj��_����H����װ��U�e:���@6��9��B"TpuAt:�i���S��a�8e-�X�GL3�����ɏR[|�-��OBd� �jG���A\�mj��+1�U/�D�˘��D�N�Dpǫ���8��}ar�/6���vS��W��w*������8������-a�*�E97IEm�#~���,E������|��3�6��6��۟��[2U�L<wr��6�W����S�֋qVҐ�īͶ���4<���>�'>iɓRcM��=��8�M4�*o�Өѷ �^�f�-I������