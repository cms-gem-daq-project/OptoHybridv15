XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7���n"�b�a��z0��|�
�[�r��Uy^�n�NK�䏟{�H�c��=��4&AZ�Mg�;C��Ȉl��x���?7����9��:��w�#�q��~u��칧��H�\�&a��Y'�� ����\z�;[��4�K��$�N��'F�&��U�c���g�8vV��Cf�|���tqgO`�����78U�tĻ���Ӷ�l
��y�A�!��I\�4t���Y~��0g)�8PȚ:�rlu�ЩL@	�'��3�&Kh._[R�q|/�-K`�We��_kr)��K��9O�F�R�76�>gn�����/\��
'��y�J�����tWQ�wWܠ�S�E��;�Г\�K�G��Q|���5j�
qX�>165�	���ar�Τ�{W�i�n��y/�3!���ِ���:vЅ(*������iF+<KK�Q���0\�~��{{8���B�~4��J�}|:�#o��a���m�:lE��EK �������hЯg�:����WtZ�l��t»���Gd仿��s�d�|W��x+��RЂ�]�&G���9�if����1.�-�&��LI&�E ��eY���U#��m�i7�o�mR$P��Em �N�G�'����	c�����2��C+��0 
V�'�;�6��7����Zq��SJ��U#���6�ʱ��Z���07,]����g�l�r�����Z�+D����M"!a[��)�n����d�]�Z�GHu����G�*~(�XlxVHYEB    4a09     920s�\���ax�L�����rxЦ���3-��(JŻ�wBĳ����=��e�O�\���^�'���̐ˠj���+g��\$������:[����=�j��K��ȑ�x��r����F��,Z���ɨ[U��7�5������g��6���w�>��7ǹ�K��+%7��y�?�Bfj��|t�x��5���͗����y� rTf����HK{u?f ���(i����"�֋�2�A�6�s�iR�Bl��H�rę�!�V+v��Z0�+�d	���gT���u�8�j��Tߌ�1ܦR�};P2 E��L�@����X���Mn�cVd�F]�η���w���O�O�HY� ��F�},��o���E���m/�>E ^�g~z�xX��|4x��<A��'569��	��������o_�?Ĭ�5S6�tCl�~{ �x�X�
.mW�X���E�&(v$�a���ΐ�Џj�y�?AA(t?dG��ݷ�"����*�i�f�Ord&��@F�*�Q�S�e�̇w����^h?F+��Uq/�c����X�`�V̪S�q��mp��	~:����.���'s�GTy:��?�-��Έ�α��6��߆W�}�i=1p� V��<�q~ߐ}8:b�2=�m(�	M�����Z
E"O�S$�ʴ���a~�1�(�?d��%�(lq% l]Ȅ|���t�+&�\6+���kT��kp�"V#���gYN�h��{�'N��`x� ��������@q5����(\�xoׄ�lK������,�%��7��5U62�{��F����������	�ٖ��l�!c,����w2~������0���|�`���B[�^mEha�	�!�M5�寨����Ⱥ�O�j\g�Ҥ��!��fz�0���Ҋ�5���}����%�B����\(B:\R��[V>�'o�p��0u��]
dBR����N-��k�����G�J#D�D�r*��p��75٦�׹Z�� �C������~��W��-�*�^��.��6��M�N��p?NrG/2�.�/�����J�}��3�3I�Lw��Ck�0ǯ���*+&�;6���0�O%#��~J�:� X�Z\�(��)�k۴R|ߢK1
�hl�˽�2N��?t���6f=�	¡ˊ�k��q�)@�J@��馚�N�;��9���Ȼ���c�k���r�<2>GH�Eo7\�
��̒>�&�-I��6�b���L��Jr�6�ķ�6�mh������L�V��,�ܤA�.�Iv��V���"B�!�u��_��7�u_���w,K!�3�Oǟ��C>�a�QI��3���v��W8�`�ʡ��L���c:+�7�e��8o'��*�Τ��9i�S��ci~yF6����Blz�f� K�'���p7҂;��e8�h�+�(_����~{R�'u8��"b�|��
�*���AK=������N���fz��[i.���CV�����*J���5�҉�T2Q�@͑�76x���}���3Y����d�9��>��О�:5�Od�k�Ч���F_P�0��=�<��ݡ�F��J��
0�����C��7T��88��4����
�
9��W�H�u��'pG�^���!��^���˷���T�g�O��Q?6'3vAk�� r�L�Hк��;�W+�)���Җr�.��q$�[ě36C3�9#��{�<�kC�i��U�-?�U3f�3�*rD.��X�N���Չ� ��@�~vi	�z�bs�ZZ:��&� Ê@�]�*����N��d���.k�rfe?o����`�g�|b�л.�%��
�o��S��Z޹���ts��΄+i��*m�ܔjE��wY��[���Pʌ��]2�J��G4��}�+�V�x��,/B����boS$sx����4$�2�Ѐ�?GN�ب�K*�� h�n��7��;vU���S�0%z�� q7�$��� �����]�
6�~2W�i�)�O���2�!�5�R�&P}�@�B���]� �.����L��b��."!�̽f	 �7�$e~����"z���6�����v�<��t?/~��Ͱ�L�ڙ`ɼ� *�C%	�vk2+���/�L���̷�+�/֜��
��
CּL��'A��:����e��3�S���2A����9@]9g��)�p�Qm�K}䰘𘽮H�{TJ��|�pB�8�_����rӠ�f5��}�r���S�O|9~��)�]]����{��8Nqw�}����	ҏA�$��u	�]���LQ�o�q�kg��L�c����Hl��r