XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z�?q�����0�� ���?��FzJ��_HY�g8���0�y7+=�>�󦓱�AƠ�:��A#^��͆S7E�߾/S���e�������fF15 ��7]�M5?`�h�#�4n="#Fꭥҽ�".��i�ԈG���ωn˝���<��k�eoeP��}j��"6拏48�R#z(��=#6x��3��l�f����A7�-xB����a=���aת�M�1R	3O�[�ۼu#BC���G�U�7�fB�|G��WkX�wq����i�X�'ۭ����;@����lD��ו��Ŷ���+��Z�Ooc��r�o!*6q��(�1A��]���}�-M`���1-�����;��5Š��}��<H����~�)F��_�@|���<k�bt���o�mr}��oH�lJ٨o�������3���o
��cN�lbn�!��:_q0�mz��?6��7B�YT�ч�����GT��VKw@��.�ϺP���s�+��$��-@�zzHo��'��`5lr�ϊr�����ƽ���>���b�p��Ӽ ��[Z�G�3�5�>,F��=�e��{�M0C��{O3��b&��������L⟁��)X���>VI�[�VO��TK	��곮a-��Dȇ��Ђ�����	�&H]%�wr|�s�A��F��\�^�3L��.\���f�� `�7�6�6��^/'߶� e���;�W���%���?#v�y8�5B^D7`Ʈ�N�<�3�Z5��(o�uY��5XlxVHYEB    6df0     b60|���hm=K���z�@���"s�<�N�57ú���CQWf�����P�u��IJ�B
�O���	�]���d���,с�3T�9'�M�ܿ:� �x��X��Y6�(mQj��fʗ_	�	�A�&r�"���e�w�14��/wމ����
6�*����n�_�����y4:��g�Q�����������!���v��V���D��Zv�o��,E��̰�@O�K�����,�%ND|��#�l�X&㏻wi0[4�o�>{R�>��P�}@ц�7�4�qnprJ���P	���H�e�ks>ڜ&�f<y��3��e*A3\��]9��.n�%��p�лF�o�<c'�גLr�+�E���{����Zp#�%Imn 7a�Ӗ]��F�פ��%�1�L�q��n{�.��B��Б�¾���3��n�{�u��*TMx�
$��;��(�3��%���8X&�r�S;�UX���X�O�}�o���?WUN���c8����s��z
����_���B|nΧ)�8Ϡ8O����j��tIF-d��1&����� �!�Q���}�6eD�L�Q�
�aX���2�U�aBe͵��\�����P�#������`	���I����\<�����^7�,v2��y����.���<T&o�!��'-�z�[ps���h"���e*�h��Z�n����Y�y�a�Z'H�$qm�T�+l�f6p�/�H~]��I�3<��*���U(v�i��oY
�S}�'` �� �J�D���Gp���كyHS�~/���Z�F$F��0�w���k_��n��b����:p�D��u�N��������8����M�N�����"�f0q<g���G��l�n1OO'�OAfI���W�ز��3�A����u��Ki�c���e�U kq8�|�uR'7&!��
��V�/�����?�0ݮR��Ǝ��NE�e(%1J� ľ+Z����f}��Cv�T^<�ꡇ{}^e+$��>�P�C7 �o�N����~�0�W�q
��D	��3[l�}b����U/���v1�����u���X�{�E\�!��9	��C��Ȭ�[���+ϖ�Pf2Xct��_���b�����S�VU�L�@V}������.2"��2j�����Cs*�2��;=���dOz��A��F��P�.z8&d��!n���\wL���7���)Z�k@&n3�����Uq)y�a�(ԍ�C@��h[L���^7جa�d������|(]`�z�\���>/�����|�n��.�I]�{\6[�SF�����2�T򚴨Nf7�D��
ըlM�=hϔR��r���LP�N�6"�0���f��[��*@ ��Ѥ}7�|kb�\������ژ���_r����ZxIo(�,ɛ8����,����-{0q٫?`|���Y��ïB���j��Sr�[mP5��Qg>duYY>|�ѳE>����A�����(��^4~o0��`��boۤ[����X����'9-���]/`Ԟ��,��N��#��Q��]��i#ަ�MyS�r�X��<��T#�u�,dI��[ۆ�T��f8��{r�Zߤ��_���~8j�%����ywk���,?���p.�&Z���2K�����,ǫ1+#L�ٌf�*�$��U\^ D�l�_w� �q� ��⊼�i%���R������-J������'=J��c:�]�T�<�N�Q`��w�(���g�m-h�q���~��� �v k �-�+���%	���Ư͔���g`?.2�'�|�H$L�w��5l�{J���Bt�����;����g�= ߃>Z�*,Ba��J�WF�� �#r�Q��q27L�|�2n[�����q�`P��t��>���aB�.�����'ne�!LX���j ��V�5��$�/#Z��#-��S.��v�[
�V�A~��֌�pۘ|��}	����n��ԕl|������Яi����t���č����x/eΣ�:�����+��m��.W�͑:�&����Ӂ��#�F����*��qwB����pvlv�
yn	g�s�Yk)瘺�C��y��٨����-�VNRԡ��g��~~�N0�U�B����\ZD��L1�!y������^�R�.:��2�4ӷ�
��|f ��ߵ�\��iqn��SW��Z�7��-�����X67ߡ�?��^E��hՂ0��J?��)K
|�]�[4�KYvо�c'N�����ɝ����\�m����L�s������;����O��4�;6�J��l�~���=$��Eʂʨ	���f����OE�Ý�-�WM���k��RNb�1�D��|� ��/C~_��U�<{��0cl�U��F��l�U�:id�^v s��d�V�����Վ�w�E�X��O#���4x<��N<�?��ͤ�Bz�s�f%�Ї��o��F��2�Z���D
���/01,�ݢ��pv�GC31t�n�<2�h(��9Ml��a�o��p㕩$��eb��K����HKvf
����j�9[��k�lk<;^`3j�������a�/�g�sd�*�=����iq���h�RdD���'��mL�.��RX�w���+���E��/]�-�t[�Hڀ	��2�>7ZZ,�l��bw���}�ύ���Q2zk�^4��ZH�e���f]$12r�X�@�#�$��
d���_�_�x�G�DS1;��{�~�WIw�@JNl���vn������DDvR�/���|f�WT�nu'-���3�Q�*�ȳ���!R�i�{TjNr�C��X�f�,�$;Y,��U�����Y�)��oҽi0A�I��M5��buc!M�