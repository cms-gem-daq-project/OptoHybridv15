XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0J��h��_9(��%�~�C��O����8��y�3�/
4��m���4#3���8�[_/��c�>�!�2!~�D�ja�o�s�rV �}a o�~�;Yݥ�hiè�|����5v꣸���?�r����%�:�^�v���R�äq�XҸ���kγ1�Y�'�����W�,�1CރSN�e��2��O���UE)[���*�v��"D*5����l3a9��]�"��[�!&w�[0���Ӈq���)�"��D=�	���B�R뷦I�L�4��O��W"�bU�!�Ӻo��-6��`XG��wY�J���V2��0Udi���dU&��QωѾ���J
�m���|QG�('������Qql��������wd	/�׹�X�?�pK���D�qv��⋧]���B�]���F"tX_]�b�x�Vޛ���G\�B��7�8YF#�ᩦ��K#�+�֏�**_��ŭ!�V�OH��I�$���\��1�����P֞����!"V,�Uƃs�o�������Y��nj%���N^�,�Teu�?�m=_)��:A�@�����H�s�b��;���C9�"ⳃ�ݼ�ʼ<>�GDN��#��IW��Z�����c�.#]�n!V��yYnx��wtg-�1v��3�-#�Q�+WN�j���W�J yW�ü�^t�K�`�vN���7������MQ4��!���UA&���:=��;������	|�_h>�j�}�c��a���>XlxVHYEB    1d51     7b0aN�ޞ�vF1]�;��{����$�7�}�o�n����E��7��uc��LI������o;�+x���N��ڄVBZ���Jl�\V�F�/�骅F�+t�`�*}����x|����ۼ"��y���g�;���?�5��7\�q�b���d�ŧt�~�$y/B��n�b�̬���.�bA�Cە�r�,��54������3�WWe�9���*Puڦ�,�Nw4��9<���'D�SC�/�˅�u�*z�`I��u����\lԊ��z������a����S(���o9�����6�|2�bD�,��3F'K��D����{F�ѸC��b��<(�U�'�%;oe��P����N�� *�JZ�~�����pF������26	����\�	�پ�M����v���K=2G��J߬��f�9ˁl�w,�V ?{���&8�7}�;԰�uq����Eg�k��v�!�֝����'��n�$�#|��`��%bT�\\��j{�hK^ZM\f蔅�t���9I� _��b<���`T�<��P��U���$c��l��7�~AAܳDۭ�uX}���+���$�2x��#������g	���c~	��h�~�pzC	�3`��)���p�v��m�6:�*�����5c��s���a�>��W�8F_�_�@���@y�]"�����)�:�REc��$�h��f�K��6s���N�N#�)����0��>i?
�#7B+RB��ŝ�7U���O)S$�3ů�\�(&�k�x�\���2q �;�Z<����EE��3�c�w��+���_�Y�^��uI,n�-l5o�Ϯ����#�e����_�������)<��o1�ߊ5]�h<�]������nBy����.JaJ������w��dw�]5�Q��U�m?,a�D6V����gl4Mp䘩4�2��q��9#n��f���e���BGp"���pe�a0��c�5]/I"�x��@�ƜQ1����M���X1�TQÜ�~G�� �n]���&E��,�w���%`���A�σY@��/�0F�]=tź%Ӊ�Hq�����k ��r��hk"򺿞X�ُ���V������fb���N��~�c�����������eoWИ9q��L��S���_�K2ϙ�Pi�H)C�K�w6��I`�ȖZQ����ս5$�ܓ@�Z3n:H�<�[�����t\��6Q�Ob�w/���4u�ׅ�] ;qDHz���#�3Oʕ�lx&'�/�$Qˁ��{�O8�S:����"���&@|�sZ'������ ����<T�>��,���͵a�o��K��r���s��ɭ'��\�*K0x��;��������2���,���1?�ŝ���!(�X��-U��W�����۫�dT�:C�zp��W�%fL%���MO���W�%)���z�N���7H�+�����đ����y�$Y���|�7�uV�Wt���9���`�؀U�/�F��E�0s2��)�OU����$R.D[@�>�}=��:��
X��}l��
L�?z?�U�� U��5�ei&��qp.'��"�)'�l�3(�dq4֋/� �"a�j�|��K���á�-Dot�X*!47����^
ݲD����/�h3�B%G��M��{s$��&rK���x��T���`��� ��a�7!�#���<�iC�}�ݵ�?��æCD�~�Sń���:Xt�V��){N����M�ʞ��<q1����U��5I'S����!`HI8�l�4yV�f����x�f����u�F&z��n�[��@�>?;�����Z��!�]����B)�L�+FE�S�_��`����9���^� ܧ�<�L�{>���^�&��T�T7���{g���K�jS3k�0_X��(b��_./��$v��Y���]K�"K�y|~��