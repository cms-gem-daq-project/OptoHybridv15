XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b[ �_i�
g}��R�\Z���c4\HO����ߏ4Q��5i�"h�Y��
w�vU�׿�PK�B.�h�%q�g���f��/D`�%g����q�s�wQM*�ǰ7Nz��M"e ЊL�E9G��+���p�um@�fb���{�ĵ��j�!XY<3�qmB�Apl ���k�B%N��жa�K	�����6���ҽ(�Sޘ�V�u0c�y���N ���+_kĵ�_/�X�_��n�߲X�&�$��=j/O-�*42d��J|��I�*�r���k�������������Ҁ��PQ�,_c7/H[:D�(���/����9yN���&�����bYyaj�?��6jW��Pj��.6�E���&rm�\����+9�A\����"�y�S�㌷�Â��k�V ���(W3�Eb�����2}|�w��;����ͬK#�E������?|�K��>Շö�,6:���/*�p\���`ܮnW`�(]�#��21|0[\0�������9�&RGgn�`��+���0��v��Xi.!l�$���wl3ga�V���?�p̣gb�%?,��C�D�h�����2@{.Y�`NWTa�����ku��D���Wﴥ	1!��0���������:1~;��ұI�JB�Vڊ�~A�Z�W^6�vߡ���/W��bL�^v�	��Q�[L+�8 �[�8_ӄ�܁|�y�S$����G�C~����j4ۯ?]X��t�LD+�*����ą��XlxVHYEB    fa00    19d0��4`bJ�U�y||..��Sɞ�Snl�Hj� p/���a,Q�+RX5��q2Fx-��w�),�#,��>y��+n��	X2~\����Kݬ�r�x��� �rc�vĖ����=���4)T�jE֞r+�����&��b����=m�#ϼ�p��o���d?78t�r!r�SԦ��e�? ���ШZS�����ք�{��YGW�����q�TMjƃ������h=���F��KA�+�NA�$xL��� /F?3x*C�^1���暸���d�o�2�a�}'�ɆpU��!��t�;���7/��Ό8�T����A�>�|/�Z�q�f����j��Wڠ�$(���1�cm�FcGG��T�=jW.���k�{K�vI�u-)�S�XgL:@�.@3�w�{�v�3�)��4(T�΄/�57�%Rls��#�dAe�#�5T��of>�n����2���dH�Hݰh�ba4Y(<^H�0���y��V#�=�Ɩ��Ƞ��_���L��b�d1����g^�=���Ѝ��j���a�w|WJ��~D�'p�PA�����@�������PK�>5��j'�ܚ���.nKX���H2��۰��'����\��ڞ���<��1Q��x|ԙ�m�����!W�1��j�2��d*v��M�JN5�_`�H��q3`�R���S�t��'�F."�?�GG��|��N���j�y���Đj��{tJ�s�\�=`���;�	�L�,)6hBg�V���җ�^g��X�L��PQ��2H����+�o]�����$�*��d� �IeԪw�e#ա
�h�3P/����R�F���^k�M�7�L�+��Y[��Z�穋�ڬ��
��,H>u�ew��nS�r_~�X����ʍDCc��І�yp�0XR:�`N�\U�{��*MD¸&�@hZ����0��E.�٦5�0*���1��Y|�"��� -�Ye�gNt?�9�Ɗf\�v'-yb9��vԕE��:�z롂u�Ҟ�BǢjs�e��e���d,*D6�"����6=y�b�˩x�
�_��8�h�:�A٥8�DWb�-�����6�
+�	�;*���,���͏��K:
8a�y���p�JX���Ė.K��@��n�*���h� �����xM%}4�5>��TN+�A]aF(.��ru�Hs��?�[co���'N
1���襽����TjY�� ��'x��F���K���OC�Ŋp6�!��|U������ �8�S%Mf_�8}�S�P�`�V$��MZs��x�C��4��Z�2�J�ZES~�<�տ�)��3nW�R��A�XN	kEW���[��J�:�C�x�F��4uw�	j�}�\����N�,	����Ƿ�w=֥�sl�zL�W|�,��,�@�5�-d�1�]��a�ԓ����,'<��ͮ��<ؕ���W��o�YC6g�_G�<��t����1s/UY��}s;��s�����n]L�\�pOw'|
1?��@X�ù�MC�w瓉�>����3U�����j���ANV�ܚBޢ/��*������Q}':<�=D�pQ~�˶]�G(��f��g��tw�Y�k�aX�U�$ՙA��� �fgueCO��V�R�>sP��PTus�f��AL������)8iaGeɘ�%M�ma�.�����n���W��Lro3�I&�q*s˭D~�GH��l�a���=���M�_���s��6/t���t=#�)��U��a�\>EO7kX�CY�1���-�&�(���J�x��n9y�yb�B��z3K� �b.��Aح`���@�!�Y�H1�aB"xjt�E�ν.7���p��?[�){x�JD�z��d㿻��}p2<.ʛ*����P>��O((*N�z�<���d���ؙi$�'�%n�5v��R�Ipc�.uP�L��H��� 0�=~��:a�Q4���K�sj��k�RE���(����ZN�Ī���O��.ۊ4?M���@��0�&��ޡE�*K�#��y�Ӗw��ø�������M~r�dD�{�K."=��.��W�,I����t���jOf��uX�� W��A��4�j9�u��~>�����|Y�c��Q7�F�a������n*�	�kloCM6v���g���l<�}��g��,F7]Oz�A4��)���Q��~��8��Ĳ;[�����p��aQ_�
y	d���d�.�_��<X��W;+��K�� �@���&��o�I	��
�}�s�ȑ«�ڒ
��My�`p/�oH�c�ˠS ���|x�'%Q�����׋u���P��۝?�	���^�ͺ�j��q�mEX<#�o/�giٖM4��-�;�h֕:�"XO���0���HȨ��|ζc�"�w��Q���3APN_Ɏ������J@�r��s52�"m:��4���������LA&+1�Fv?�s���4W%��5*�t�L��ɏm���*�-�ާyA`g�ѹ�ʨ�K�*p�!�	Pr+��2G�LT5E�e��:'��J����j}���47幺��*��d��~�)�k����M���mf�J����_T���Y�,��'�]'+�,7����-�K�n�vj!y*��y<�ʯ3�szW��~&��>�ܛ���a>�G�c��LX�v�Τ6�wm����
���Cá�4.7Xv۽rUXc�ؤ�����-Q��&������I�+3����膫��)���6M��t��Ѹ���/�Nb�[,����t���z��W���d@C���D�§W�����;HDQJ��7��2*���� ��g-��K�G�+��[�tr��r�ؘ_�d���8�5�C��]f	��j��"�b��ĦAj�=�I5y�9{��&���O/���
=��nT�����پ�Xq�P%j��S�G���(t�z�7�3I�}o��C�11���g��<�@��h�����h����"�h].?lW���Kh��/�\��T��.vU���H�|����F�	�-R���0/����Qĉ�c
�4B�v�S�b��gh�~v6��B�B"����Ѳ�@G�̲��Y.�?��)��3�ǀ�Jǀx�w����B9�F�����4g�v� ���I54��-anyv}�a���9@T_hp��$�:�nq���lO=�֩�%g�ag���gf��:ry/�x#l�f��B�7_DO�g�Fsl�@�4�|G���k����H�!�8Z�"����*�c��T��(f*}�u�}�zn�U�+�M�.2�ݻ�]���+ZJ���8����X!��<"29;���+�p*x��WO�vT6������:���j����B����gsY�1鵙�\�*c�krx_p0E8�(�ù���ӡ�;�AB����%�"���į)�&��1;�D�^��;v�o�E��k��/ǑP\C�k�x�"Vx�}\j�%��v#��j#��Q���˙J�7C�bY����/c�):d1����3E�в�!�gQȡP����N��b�������YF[�������k��M����y޹«��S��3@B�����{A9w�j��rx�i	��!j	��ѷP>�e Ut���p����=��$ԺU-9��N=DѦ��m8슙cɳ�W"�_�3dN�)s�I��73<��fDB.��9�JGb��,��Ha�CxÖ�ch.����⺢���oϥ���iU5���y(Cg�[i�C�t�W�'�9��y�%߈K�������5��Y�ې𫢾tA�Q5tQ+>�^���ڳ�КE�Q�ST9�1����봊���I]�1�C�*b9�d���	�|������;�+&[#J�T��˵4�q��I��BR�I�c�I�T���n�d��?�a��vq�qO�0T�˯;+��d'�&@�9=��y�0.yR#�Q�$d?�1��q;u�J���l�.3ҢП�!�ӳ�*�a	����F�a��Ӫ8!�M���):���MO�c 0g�ǚo�N�;�}-?5���/�+������i+�ZkW�Y��1���k���(ȇ�5~#���|���`_�߻�rRŶԈ��ytQJ�w�<�iW�˥D�7>�G�M2e�m�P��hf!�ŤT)���n���kC���20�.\�  �ǵiR����78�R��mG��u��Y�.� N�*%Ay�E�؄@��J�'	�X?G4��������l�ϣ'�?J9�a�]P)K��;u�+^d�k�_�Fg���8Eʈ(�EX��Z����S�2��|�ȃI ����s��j^6n��ǧ��aA�7dE���������r���W=��a��T4�f
<���d.Xb�0�bg��ˋ8N��\��'���o�Y+#��AsX[:j���Q"�ޤ�p�r��z��U�V�|�a��R$��i���Kiy��êF�3|l <�&��RME��I)�@�����O�^|����t@!�`�γ���Z� �\��?�S���)�ڡ��igR��l��ODCj��z�f5�7�蓶�n
+Y�b�!)�Z׻i��e�l	0i���q��*aRl��A�q_.�	�6��HN��X/�	t�.�D�uuh�x�u��"K�O#S>@�@G;�s�#~OW6��&���T���9
טm�xO�R�V��������	Z?��$���V�Ȣ�ݹi�re��Ȕut^"/�Ou�,����Vg���*��[�N�e��=�BӢ�!�n�Z��(��
���2��Zu�B�4���<ce�%)z��7D�@�t������ۉ|�U��2Y�ە��Ϗ���'__2lK.<r:��)�$�4K�dS�B�M�f�����"c1Z>쵒}�p��pQ�L/����i,��ӇZ�{���}�o���q=�I����ޓ�3�5��?�a
3��H�𵮼�%�$+ِ�xN�_Z����G{���X�x�����1�(/�.⼏�m�x@�������������3k��6n?|���1<�������KV����@m�Q���%gO�{K9�Bݴ�w�\q˖�`E?�aqïtՠ>h!k���/��N�wDOif�ٕ)-;c�^��e�S�9߀f`L��X��Mܓ�	�k�MX�iD".	mM���I��$�����X7�PE3��{��T!st� f���a��,��sUr&"�t��镭�j/���4�I��j�?`�2�2���}�k^�ޠ��C�F]A���n{��ڡ�%G �9�|�W�?�HT��&�,�hku�����-l����� I�����l�hu�}=�"��R"� T)�� ����NmD��/C"�3���l��rȦ�t\�;�� <��V��q��Zo�iS���xe1��^Օ��iz��ו���+Uˁ���+u勵�M}�]���V̺�b�d�Jf+�o%��b��.{�� ����w�&Ί�j����f����Ш�*�s(�r�8�ia���q��r(�<�����<�\�<������	!����I$����rH��y���B�%Q9&�����-D�q���<���YA�Z*�W�ւ@ ��DJA��k�b���<�A�0��2��iC�g�q�?���0�]<R=�r|��Bh��(��^��M��26����=�Ʌ��π�m	�d<� $�E�e�|G#��i�"!2'�v�qM�8z�}�m���.6R��'#�{�<�q�� �B"�������]���@^����9J�F/: ����C�v�$�Oĉ�Z� |�U8#q(�4�̕1���Jx�jr��O?F���k�vD�뚾��ܮ�{�:n�\�L�+�z���T'ֆݣ�W���V�5�@w��N��k�&ܵ�#՛�ࢩ�0w�a�hq^^dD��6��y䥻��zvՏn"R�}/���v�U�q��m��{�.�v嘯N�;�Nv|<Ű��H ��<�CU��l��>�a����嬘I7а�37��'��Z1�q)�������QN}��툞$L�q@�f��V��eT��u�G �X4�6J����������L�w�̎X��/N��<���������w�����.�w�wŞ��e~cqE�q�0�P�����k'�{/�nG%�p��]ټ5����ƩeB*?tJ����Z2/*q�G���O��S��0�~����� �"��O��'iB�Zp\���z�Ǔ�Z�b8F�#���O%��㘋B�˨�a�$�L~��?�S�(A_�{v*_��V�1���W�q�"'o{T�h�xn&�j�r@�Y����)��/ B�]���Y~C�������E���ym�h�x�1;��阩�q6�l���ŵ� ���H���e���Q��W$k�à-�� /:�Q�	xe��;}̉D�;y:l�^LK�]e3�̢}��ڷ-��@�8'޶�B�k�'؝��A�k��Ng�դ�ڐ�1{8ɫ��{�:��H�;XlxVHYEB    fa00    1630�"���!�&�и�PX��ᯢ���0>����Շ��R.1�i:Oƌ�Cj-�b7�9�1띍fp!+��n[��0@�v���=M�p9OD���!uȌ��H�����bi)t ���a�2�N��0�PB�� ]�����G�{����.�Z����y�$�df׹o��� ^�c4�tn񻮾��qX8h�%N�n���a�zP�D�w�W��		p�&9��'�������~K���l��%��~r�h!�W~�?��$�љ���H��5���㾝���/O`��O���G�2�P`LUIm֥�C:+y����;�T+����y��1�2Q�p��������01�:Mxn��r,P%�9RB�q"d� �0�����4�� #HI��#F��/��s�t�ƴ>J�AG�88{'������[?0n����)gG���z�È`"0�lGt;}N�Em������c�!p�.���:k{`�dG]��v�� �h�^i��r�衝i�pq\Jx��Y����<e�r�� R\  BoY����h����6b�<7u�����-qq�CX�%��󍐕��)�k��J���#�PC��w����}Y��B���U*"�E�_&I��R��#\.^D|����>nL�j%�TP��^o��f?D5H�dDm͞�3Zg��G�g��VYd�8U�T!v$�Ek�7���g?1hm��{Ό@HCx@P|�#s���8|�. ��h�>(br&��A��t\Ƽ�o�RQ63k&-'|�:��P=��4��%6�}Hz�y��o�{�v'l��r`��g�*@��P��A{V�D�M��>M��\�7���\@ݭ�����+��a�#"�F�祝�5�X� �����Ul���X*�K%ϻe�,�Gz>�]��'��[�J�)u�������6�@ɣ)�XV�'��a�y��	Wޅo$���tp!�e?�U#�qyZ,��b�I-�<R�n����J�t^Z$�dp֝�����}�ܼ����z~��ۍ��ʁ�h��C�+h��6p33ê����CZF/�)�ߣ��*G�o��n&����!g ag���s۶-���*�С����1[P���	ƒ��'[��'z%
���ni���+�Q9j���D\�B�g�)~�MD�^�.m6(yt[�jOPS��#rO8NF��7ι`ޤ`*�?��[�J
�5�'-�s�6������ܯc�``��F��N�sD3�l�?$hq�#��<�2��i�U���7��iQ��Ȳj��4�#ZLɨ8�f�7��*�c�u�~+Dy�
M`똫[m��ٷ�eBhpHCS�
D��뎀�W���DF��N<y���R�l�b�	���3�/�u�1�&�R%�qdJ��wP���{�`ʚ93-�XW;t.��	,��C���&�+,Vj�4�%�0�b!��F"���geKD�i�#9�[.r�_8G�w_w�8�H��G�pp���y[�1	�:��,�C!8;V�6�g-vJ1e�g>0�@�%g*���^�Qc-�^��K�^z�}�R��J�޺��[�������b� JprĔφ8
�5{3S��^pWw[	[��l"+�k��jU�7Gx
K������=���ݍ*�E��Q����������z�����Ԝ+��MV\�*��%�;���e�{
k:��(��Y��Z���'�ߤ��p'��/i	��{���'�XWy�<����yAd"������s"�c�mn�! �=L�I�� �|N R���Jj��n@�:B���f�M��9C�6k����|�9T��,h��e<p����M�^:�9�"����ae�1H�p<��K�W;���h��a4.d/� Ȏ���2�@��"-���&,�T�5�p����*�`�8�`�*ܟ?����T�$�8�Û/�I	I4[]�pw��pE�(S�VGU�G�z�����'a�$��ㄗ�ąP��:�Q��Gw9�{e9-�)���!|L�z��k�D�fa�G�=BH��6��s�ڧO0�ǟ/���gF'`�e}Y��iM�PԚK�����k=[Z�7 ��v�r������S�@�,FGP�i��,WE5��� �@��(�O?��V��s/�D�;X�*;��~y����ua��Z/�� Ɏ�"�#Gs�@ %l�]b�붷����D��*h0[!8XBۮ.2�ѻH�l�Nt��"YDKE�'��MbA���� AP��4�G�����q�K��D�Pd��&���������j��+�1�z'{�as�`	�,۫�<��7},Ă����ǜ{�y�bF�4��r����T��a�l��� ��ύ��#jn���fK�$�I�7����*�����j�!���+�l��a��z#��T�y�Uܕ�6[zH�C�.�{`�_�ICs���i�.$?��l� ���'~)٨ �0�"W~�$g�#�Bdf��^���nIPu��G������S����|��(齛����%
?=�wLχ2��|*����iǶYn��EHH��O��+�o�u�d}?_��;����y���fT�V���������Bز���^z�n >u�M>�::	�	E��&��Nش�D�a�h7z��17��{���Ĺ[˶�9���F�����WlC�
u�Ǐ�32�1r ܗA`�Jӏ_j��m �۸���ք���-"D�;�M��aI���L)=���,1#��T�����?��&NM�ↀ ���4�.�ZI���Y��<	�L��>|"�1��pG1�C�$�C�ϝ�"�wO,�;2?��t��j�aF���Õ�����N�-�0�Ĕ��_��y���U�O|�6>�T�=}P9��D��l,Z�Z%�-��҂;����iu��o7|��{Z�5�7"<�ɖNV*�Ǯ\�*s�/Vs�C@a�u�&/tb@�e�bF��)7m{�107q��U���M}q��.�&n=�C� ��o�I)c�ys��*į�)�[���Q���B1<I�_�`X����pg֊����UF���-�	��s��:;��{X�3��^=�+0�\"�u�ʙJ��!S��2��f�D�������L<��c�as'~��)��vm�s��Ks�;b�������T�ӡCryqb�k���Y����~�5!�R�C�pb~�& ���n����G.�޹C�Ň`p�Վ�_�ok�d��� !\�}c	d����ZU��ᬸ�r6���'+[��ah���;�+1��C�1}_����WFg?�Y�/�!�xPi���;O��L��|w��XRt�~lEx��k3+�]��WqV����������/���8��Lm U�i�K#|c�|�^W�C�N$p�������?j�[����_A��ɠ��t}�G T�Y"{�C�*��`���y5�;�9�a�x���*/�E�mI�]�����uL��u���4?
��k7
�Kc��̗��4��JeC�	��QS�x���,
.;�������͞��V�EǘĈHS� <��%�כ���OK����'}�Y�Áț����n�= xP�,z�5ʹ�~���#f���7���#�6�Hv�y~��/�|���]��v��}��W�6I�"+˨�c�ԾK�������<�_c�]�pZʱ�ϥ m���a�ǂn�b�ц�8�:��O�Ԑ�	C�Ra�d���V.Z��1;U<2�SvJ�^���6����d��i��7b4�H�㻷�T��~�Sf�n*��������U���J�gZ�&��oY��5���B?Dw�s;�&X,����_����P����V��K�U6p&OF����S��~��ݡ�hvk�����9){��l�O��Y�X���:} s�q� ����*�&$�h�,.ⷡ����n��P�<�� s����f�C�D�z�d��b��7����(�Dw�Ѝfܷ��Q_=Lɇ�l���g�>g����Z"t����>F�ѐ��E!�:��ooߟI�œ�*�A+}P�n��]��|t�		u<>�=	�5=Ŏe�;��	�:j��Tu�$pjqs����1�$��������6C5+�^5��[�'2�<��Ί�Mf-��ܬ�T\?lx��ǋb�`52��T�U���9N:����WBt�ʪN���p�L���
Qj62,��΢J�.wR��B:6nNYl�����R��2�=����Hh�7��.�^ǀ���ט�4��#�)�Ɨ�0�����|v�Lm7�����������N�M��A��'R�l{�4h����-}���L!�V�K��|�C�����U9FY�i	)>���Z@**�Ya�w�N���9PALm��\7t��\Rc���:Ldu<%F���!�~/��bB����q���巹�� N��^���1���X�(G��C6��p� O��R��&T���CSo����k�E9s�Gq��_��"��ov�Rb��C���Yl)j=����N�4͍���;��_�D�k�&u�3�� �q
�OF#�,��[3@��U���KS�����G��>�b$a�N@�p�ǿ����xŶ��J�:2���&詯���2��2f\�4�iH@�
��=��)��������)�8։��5_�NkD!w�o����������"�,4����պ��,�(\^Ɲ �D)-r_��]���i��=o1�hW|w�W�Px�>���:�,�ζ���.�?��]��5�8 VB��繻�8͋�^=!& ��.X\Mn�_��v*ǅ�E,�#���1t��N�����I�S+��Y�Qenr#$�߅���1�l9�]D�Ѩ��dk�X��}.��Vn���]�ᾌW�p�j��O"��G'�S�^��ۘ�դ3UC_�]Q�k��\H�����d���l.��{m����\uj�I��rU��I��J���=�]jd ��N�.�بUC�����-̴�z�`�ߤv&��u�i�&�����9VI�z(^�3�K�AF��%!���j�֍��&ӟg�|�s��l{�i'����[ۗ�؎9+&�j-��:����5C�M���sƳ��ѻ�'mCP9�Y8�.WB�16��um�
����#�B���52U#Kk��,jz��xO�x g��@O�vG��O�D�݊�[h��d!\?t� �����2�Ӡ&L>:;�]r�*��f��0�ډ��8d��c��[��K(=�g0 E��v�w>�j��
p6����2��͏"�dy8�βlϺP>�,/	y�m���@͂�'�M���HA�̣2=դ�7���+�E���H�#>o^헯�O���2�YV 2��yt��
��)cUh��*]+2�ѐ\��VSr7@���ȒyE&��s+5؅��Dg�Plx?�l�X�$ ���5�XsT�w�t��7REyx�1�v���-4�N)>��O�㉚�Z��?GS�ǂ|���E�od��0r����|�nM���A�3f����Gu�}�'�M|�U�n1>�~r�!���y5�҉_f���ʼ��gp|O4|,:�q�zQ/~�*���rW$��JIΔƹl�m&�Å����|�-u~&L���˶r�k[_Z�+&�3[O��x�Z|��C����#�pXlxVHYEB    fa00    16a0ea4��"F'�y��G
�S�J4��PL�7�a�
y���Uj-�����PO�SYQ�z�hF��$�&�v�%�[�6�{NP�|��Aʐ	>�R��(����|�Z�/vYˠ��s��)u��� -�b��F���VQ_P��Y�@�;����']��\�A+���y���ot�g5�m�j?�_���E�@?��r�C~�?b��6�"wg�U.�=������v�h�H��QHTY����
�Fކ�}/���)GS,�&��dۃ�$���:�$Oñ�7b�<A��V(���O��S�L�|�ǟu��u�mK�T���5�L �.q�4��#ڧ�!=�H�cn‛�n����pnT(���0;!d0���B$�!�?��ս�;Pi�D���`Q���a�s��@Ă�Z���ܧ�>����cBoSۤ�L⚉�����:�{���m�뽯��#��A���&��R��jv�'��7�b�����N�G5?�ץ�����\�<��֘	���`������o����*��[ҥ({�<?����/���؀�c!vv�#�F2���,�<o�8y�.i�\�Z�%bq��F��'n���j���'c$�n�n���L���6�D�A�]��C��I**{@�:��?�h���G60>��l�a��ީ_�u<vz���{�,"4���r�<���S�h��%(ǉ���+_�T��~��e
F!������[�'s�U��%.r��ު�R�E�Ͷ/v��/���\�SNP��Cm�.�|�\h�!��۔�ꜙZ�����o�y
�bq�lА�Ѿ���'��xL1���M�h��/C�c*P���af�;Q%u���}Z�*3��/�@�>��_/���]����n0��[�1F���� ���$�z�G*�����7�*�Q�Ɍ8�6�\��~��?�@:�jt˓ek%f"�TJD�l�e�C��I4y���S����Q�_�B8XǬy���J�9�,3�I���/�-���U��Ҥ�+�c��U���to����{���0Z��:W��N��犄"0��>跇t�fIW.\̕5ׂfx��;pg�,jm�:�Ȝ�]��� �L���ʣX	N'A�^'tDްz�mM�r�
�(t�O�c�{ӵ�rB	H`��9��Y kg�DI��t�3�W��Me��M��G3�\k�̯�A1��e\��l�p�gou������X�Ӿ��EeHO�����.Q�i��Lݐ5�g%ݚq���Z��J�0Y�W�µ��|΄R���E��[�L�M�$qZ�f���J���*����]��&o*Y�Y�G%��kUYƷ'�����z�hSt��!z�7$o�I�T��5I��t˩	��qg�Ru��3�����_�폋A0W���BZ��&NC�\:�@���Y�f�v/E�Ϩ��	���}7�u���Q ��ȥ]x)E�ZlN�Qr>D�0�{o�ߺyN��{J��L��x�-_����[1�`��"�m����ȱ0i�@�n���ꋦb�t��m��m/ݛ��[zS)�T���B���	��m��y�d�?XsEz��@uSU���#lo�����vqa�\�,��	���� �?|��];7�ke�}��;x���l��3�h����I[&���v�������jֵBg"q���R^,w�Wi��ީ�/P��W���L2��<�G��Ő���{�ҍ}�d܁�c���|:-Rt�8��#�������(���ІP��l�����И�rH�\�uC�8'N��ٕy�ԟ�i�$�"�4G�4.hC�(�|����\��+��0o����G�ü��/�'Tͫy�8Q�U�(K�>�c��d���<�.V��*���R��]��7K���èL�Y�c]V�8,<��O�5m�W�P>s3�L���6��� �M`��e4�����D^>��#Jj�+9���ĝ�7�h���n{��/�p8���~i�l9GS~iZ6��.0һ���=!�#^���7cj7���P-��k
Pv�Oݝ&䋅we����g5cc
���	����Q��z �Gx'm�dmcJ�-�>6*� �M�Fc��60��+��i���;.�e=n��n�(�� uR��������=�Z�7���kツh����j�ԋ��<}����b=���M��E�"��~D�N	�e7Ѥ��8wcj ��zJ��j��l����ݨ��>�ƾc:�	T�Rj���A�D+��֙IsV�|O��5���2_b�I��p�)�_��!g�߆T��1\�Ʈk$ToF�JOaH<�89�)BB��v�3��E&6軖�]qg� ~G%�k��+Yu��YQ٨�r7�L��K��V����&
L��� 7�aO�U��SG�e|zt:y7�J�T�x�i�R� 1�����اf7��`6�E��D���ý��:/J_�?a�❑Dc�l�����ްm��?�!� �T5��7�|JY:,坫�x���U:|�VA��|��,l^S�:θ~x6"g�>L�jdd�g?ة��]�r���5^{�aR2%���f�YI'w�W3j�w'����ނE���5�f���K��Ǭ4VY�ߐ^�Y�Az��~��v��%������O����f̦Z���^�d�.v���S��D�����I`�X?o)��4d�~Bo-~$/�D|X�<0\.6�����Y��K�X����95.�j8g�2�M�-��Ih�?"���fI1J�5W�"� �����k��Lb�S$�,��^����x��,^�oI}B6��e�7D�$��S�	t�s�������Q�����/���2�{�0k�iy�?�!Suq�)�;���,��<#@�ϧO7�2I�K{K��?i�T��U:�Ns�}�������H���?_�hcB=�#�a����H�鵹[8$��[_�K5�:����FS ��h��6U���sp��w:=�6Q۳�RȐL����;{�Zh��u�\�LI<G��s|IǙ���5,���.�n0������L���F��4s[��ȳ��ñ#	K��y?���O6��<i���� m5χ�"XU����=.Pv��i�u�|ꎮ����Tue��'?�&0Ѷ?i�ܣ��P�9��56u;tЍ���A�D#���c�Ҭ��0��G�U$��h�����7�*�N���TR�����+s�h��'?�i͒C�)��~h:���4�kD;r�9��M�J� �kA<~ :+vb��S�RT��b��gr����))�r�E�d[a9m�3:��{V�C�mljD�����B+�Es�H����/,�ʸ\���N��(�������a�����K�|5y��ތ3U#g�ƪ���ϙ��$q��^�˥mo��t%�"7Q���Lk�d�� ��Ёoؾ�6`aD��z����Q����N�Ӄ� �ig��Tvk�~�N�X�i�.'��ƃ�>���� �JZPc%'ts�1"Zb�c0չs:'ak�h<v�&������ax����A�D�J�c�cD%��b���{���P�f@ԛ��^S��Ys)yn#"�&FW�S�7\���#�$�7;M�������c�13^�Ҟ�I	�'�Z�=	���ȍ�W{g��a�8i4��c����)T�·��}i�gɝ$:�+`S�ӝW��
����5�J�So�ii���/��ȍcJ0�2��@o�|~�8�5n��s��@G�tq]#���ӋsjG��P��.��
F�?B�N�
̯�Mw�����r�>��|�:ia�i2S�I��TZ#B�E�wW�k46:�%�i�?��X��5�LYqh$�v��u�V�]���Ɣ��2���2R<�����w��#J�ۈL-���7��v���?(�pȋ7�_M#���d7��ٯҩ�x�s�C���{����3i�A�ƛG~��pN���G���Y�$*��^�ǋ�.Ə��?%�gp8�����o�s���Y��z�wdg�N6z4<��N�(�IVz�+�~����FW�Z����ﴯq��E��a{���z��ѐ�@M���ԓ����s�4;�W��cqf���/��{F��A�%n����A�$��p	� \�o{9����x�Q��bt�g�|��qV	}P?Q<��I�EX�������0��1�ֽ�����I--��D�n8�áT%	�Po�OL��?7m����*�&S9���̷(�o�q!-_����5آ����������A�f���8N/���_'�w�v���N���;��ex��)���
���(ߺ�=kf�B��U��ԉ���L�LV �?�EF����yvS~�Ǫ@W�Ď���0�'����x)��3�2�g �9L|#,='E|Ș�!�8�(����
]��W�ǯkl����� ��;YJ�k��w�(���(AG��LEG�oR7��9Y��e7]��D:��#�V$�e̗LB{��(�ƶ3�Ry}W*�}���Y�wcw��+FI��ɴ�P�+�sA�4���H��-Op5��칈ي�9�������Rnk� �bo+�K]AUWғs�ZE�(n�h3����ޤQ��"�Sg�|�=n��x��s�[)��.�*-�0ܹګ&4R��;�G͖	)��O�:%u0.�S�7o,[�x��6�,x?V3�h ^����\�����8������^8[���x\XH��+Wڟt �g
k�Y$ȱ*��/,��Fb���7�Q7��y·���
`�����5a��{7�m��Y��iE��ޜƱ�� ����z,Yo�a1p�bc�_;Jgn��cז$C!��]M~�������̐���'�"Lo-�E�Zפ����D�j	�U3�B�p���t:Vm����y��[�t�6%
�����l�r�GXs���H��y�����������H ��&	��6�U�嗹�5���.j9�����Tt�B��#��	��Tx< ��tL=��?�hD_R1*�)�c#�M�vX9y-����f�Pw��9��dG�"�m��ZR���6�w�:��t�j����	<[u(q���$|�\��V��M��	@��~HG���G�N� ���Ɩ������3�� kxY7��l��-��y��j/ͨ�nn�>���pnw�9L�؛��KyRh�)cC�4N+�3:�y����	le �	d��~+��f�*viQ�ՍL���=F��ꭵU2�9�t�	�r�0�K��Kl���iA�F�lOi ���H��qÚ�ԝ���Ev7�ٗݪ�Y �sw��?]��T"��`�$�p�4��2�9l�/@��<nAIz�<za�\��� W(+ɢ兑ԭ�8�0����ى8�$*�tj��Ӣ�`�����}�f\��+���ϗW�~P� ��H�zc#��ߐK>�dа��Ҷ.�������]$��wWûn�8��-����^�'��117E��	i'ȧ���P�r��� �0�|O�WMՖv�L�1ʂ�����eD����*�e:�	��qv��K���|��=�L�T���fq�zM$s� ,�D��S-�lg�@C����C��}���������.]�a�g���v��8�&���Z�m��y�A��VI��Z����aC(Z O팠�ܒ�#�"|�s���82��XlxVHYEB    2889     400g���+�n/������匋��0�[8����w�.���F�Q}�>�m�O|� (H?*B� ��M�<� {�� �1~��N@�D��>����u�S�f���]�.�pƂF�̮�'��C6F��R�̍$��}���ޝX��*�g]�$月����z�d6� KL^(�D���>���,M�;�,�<'��3O��w�ˤ�+a�u��a��X[�����Rq�����0���͈ b4�U����Y�t�˱,��I�g��.�@�=w���{(U,�Q}�� �3kml
�(9�E_o�L]���8��>�{ ���O,��ժ�d ��t���.@`�t	}i�5��� ��r��J�?դ>
Q��0��~+��؟, �?�dhg����0����8������rq�3�+� G��u�_ E~JW�dj����
z�w��sM���p�k��=���1��P���o_� �$e��!=c�A᧥���S�eů������c���{��>�q�/����p�;�c�4�4���vEU	���E?g~����-��&m��k�}_���w���el�X�a~�8m�#Y���?SCT����B,L��T�s��a�B?)e��J_9+� z�+7�>��{�U�a�����~k6�4��$�Q�.�8C0n$v?Mi���!H��+�Mx�ގU5#����<�z�=����]&��[��5Yڥ��^Pέ$��3��[�`і��yi����tU�e�d$ʆ萢#��X��� �PX;�du�D�B�s���g!���Yc&>"�C��]��4�:b�ꈂ<)g���l�'Z����;�!.M'"!x8��jjGܖs�/��Ў�V��Z����Q��t	�g�C��mx�3s,�`_��IN�� ����N�Fhh�#~��r��?\
�2Ԣ�w��{7D<��9_R��o��g�(�ަ׮��畚?hu��y"��!@	1�_['`�b�!^m��_��[י���`�E�L��Օ��N(��