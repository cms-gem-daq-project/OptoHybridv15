XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#e���xO�$ٝӗ�O��B E�}�ã9�������4}����8��l��-r��y�< d�6����z�V��O���u�x	#�.�Sy���J74BXoA�K�(����_:�Ӏ5
��\�7c�Q���rjq+���N�3d�Wuȗ!hr��<�J�<r��D���Qb΂���`o]��;��U�2����E<(tn��ܞ����D~�Gm%�:7�I��u/pw�����N�0zB�o���	?�K�j5N�';��v��ji	�H�>n_ɋn�4#/����g;:��r2!����S�2P:�Xۅ|��"���u/bkM/��c[Jjf��Bי$*�l��\p���]�"݇)Ǯ�C��ԅc�����[u�����/�M��A���#!! M抢�(w��hA{�+��M��97s7��1K�ezu�#G�*`& ��_��]�l��s�ZEb%u�7K1�s
+-S��'�B�A^fo���l��m�|�}Y��:QLn](կ+����iΪ`��PW���MP�^�DPKk��T>��ڹ{���}���9S�X
��R�a��r�Pڦ����e](P�>�6̰���E �����<Jr ypY�j�K"��o�S]\?�ca�^ �����������W[Uo�R�d��5D���w����h*m�Z�Þx@�0����g�<���%~�y��E,��=�X�t�˩x���h6�������Ӓ%�#�Kq���X}j3� �G�XlxVHYEB    1041     4a0���ŝKd���-����8^Ɖ	���it��3o�:m����b*����IA��=��ҿt��Deb��!{� h=�n%���q'�� ��2�(��H�_gY����k���f���T�q05�Y��/4������|�"8�=�݁ɘ��hq�H���oD9l�Լ�6��O00��,R�s���G�`1�E��ލ�iҋ�xߧx�K�7f����ڥ#�c.t0�շ�o+xs�쁟QK���B��p�]n,t^_=�߾��ս��x>�  ͷܽbF��[_�f#?tr��t��;.j�k��#������7��(l�"��[��ڊk����\�¡�q��R9L.j�'�Xc��ci,�Xo|��Ϋ��n�V�/��f�>h�]�(��p��d��a���K7��S�W�)���)�An�BNf�;J?��Fb#R���P��_q;���}u�~~Y��;L�-9�����/b��(�>	��1��a����w�u�V�̙&�bq�i�٦�꩖�"(&A�G� 
g�bE:GRN����-o���-���u�b����������g�Ս�YO���|D�`s-G!�ץ����wooj����x*� 9���~��C�>&���������v�R��~4�ęI��ޜ�� �g�1�p-��k�6���|;�k؋��Jy�E����t*��-�*��%����d7 y�䗼{��(�l��l������P$�T�+n���~蜿������`��ë��q�	�Y۝�)��:��|��J�l-/��e�ճZ�F %>��#w��Ky[��;�p{�E+����X�_�n7�*�; z~U��c�zb�Q�.�n�ǚ�U�u���+���?�K&�Ѹ��F嗔 g�\7�Yud����:ST|��@�=�:����Y���~�߹��l����n�'
�U���-��0��K��f�bN$��8���Ԩ�jl�N�A�;�����~4����k[p�y�7L��[��#k-~m�ig�$��5
���ڄ#~����0��	�`�)��uz��/z�u�?߫3���4�2(�,�~��Ų�(�8]t�D��&B�>I㩭ۗ��KE!wET�n�d�5�W�����|i��]�O��9t�x��+�;�;��*`�i