XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������$U�k<�N���dY�7��.}"�m�u܎��*�ǎݮ��Up���r�CP��ّۧ:��6D�v��|���n.�[>�)t��F����S��>PI�*2<��r��a����-א#.r�]��\�So��v��|ZzX�wL:#��	MAu�6�w��t�ٗ���<G���������-l�0Od�^����Z�%�3(��
�k����ːH�~�>���:�CAU�e?�œ�Lk��%��ٚ�d2[4E�l��O�h~���%�o-��:�}Ÿ�C�nc�f�#��>���Y��O���بV�7���ԟi&� �dW��>�K4�P�-½�7�p�˫됸�����Z+nekL�fT���Y����Jȳ
e��"��G�U�>��r�nX?E���p<	,�z��[K���-�L��)�j��ڮ�O)e��<�.uf��ר˥�!<V<��ʖs�|r�@ц"�5H�ط��޳�5����M��N5�F�)/`[����	�q�
D��UF�0�dͤ�A&�Ꟛe���z{�@FU�l6B|QNo$��4��Nt�F��}N�!�,����!�v>]���ѻ3J���H��U�a�@��BG�b�y��m~��yt۲{�`��e�����y��K��j
��Զ��%�]��1(�)�0T� �`�T4��
��h<g�r��ٝ��'�h���}���gL��pIl�����qsE`l������b}�-�&���W;
���X>�s�z��SC�oXlxVHYEB    156c     590'9'F�V#b5�%
��|�DsA�R�S=�ݥ�i~@Ԃ��H���}�z����Tޛ󢥽�w�$�T�'���Z�ڜV_���i|wh�.s��/3��Ȋ���j�!�	�@��Cs{�e�~�3�n$��{Z����G�K���F����X�)k�(�%��fR�P�&Qo���s	8���?$-�2��K� �<i�qh�4s��(�7U�)���v�w �N�]&�(�����T8��L�˄΋r�$��v4��H�,F~�M�7 �c��,\���}��9�Zr� �H@
U���6�[�.���o�I��_���P��k�5�hey��4��7����i7�����%�d������t��Ǳ����b�v����������o؄D�_씿Ö�}���:��� x���J!.��:e� ����������aZ 迠���H�1��ƍە�˖Z</�Z,�Mg���;}�j�����D¥Hh���Y��P��P����_��u����=й��)#Z�]_�?p$�T!���{5�_�kP���.�@@�ٛ�|z$�T#qS���:�~�m�h�?������!��R.��3���=~�ţ%�J��yfkV��p�մ7�<pu��<@D��&����{*r���;�:�y���<�[0� ��Gs��YR"�6;�JoԱ��ϲ�[v����;+e�<���+n������:-&���.�\][���m��� ͙0_X댝8�f{�C�C�dr<�q�r���/|ӧ�f���z��ʂ���%Ps|��]y�H�h0Ⱥ�/YCֆ�ۛ�_��MHڞ�8�di* 4KZr�,����p�(�:��j��廲�+��oq��"�2&�������㻿�9k��S0�ن��z�I9��-H�G�\6Ew���ι��|X���`�����^�}�+c��~
�gVBr5���#���p�u�^;V�L�:����%1�f����j@��%O����{5�};#�0�B_E���#T�Qn�܆�b[ȷ�����6|bn�E��r��P�s�+3^
}r��j�
���"�{i�w?4qM!������iTn鋖�
����ҊB'1&,`Oa/½�ޫ�=ǂ5������^�$T�g+���#�;F�.��w�;h�n�ݾxWk���e�rޟT�÷h�[�m|ؠ����,�1%����Pp)�����;��k:r�G���o�8CWi,6�3���ظF--Q1E�3�����at��/�ȫ���ۯ�_��Cy9�Q�������S��ٳ,����o9
�yT�.Gq����U�`a����� #F\S���i� �P`�l߀��wRQN_L��l^7�);T>M@I����.�