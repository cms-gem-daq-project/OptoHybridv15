XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��pV@�L3q�D"a���D�b�FUb�̅4<�����Y�8;��k4:��6T�����'�\P��\w�+Ln�I�0��6�9�1۱]���q��N9S�Ҳ�v�u�St�7��S��Cҋ�V�{m�#;��~=w�W.wa�9�:�uԺ:0Z	q�ĺf.��P�L���O�lJZ��/�;���ُ�A�#������#ch�s�����`��̘�E�]�E\��C(��v�6��W��悈�ԕݒ��(ōY�g�Ճa�����Fp0���<(�ʒ{o�]���.<���V��V&���6 /U�F����%��gz_��ѹ<xIUv������fj������ʈu�7<������i���_��%����"B�]07'��S�yCc���S�k�N8o{�h�<�&`^�d�nLt�.jUBt�#4Z�łt�Ĳ�U��,�r�?���3,$��XblX�A�.�f4TƝ�GkS����c�v6�U�J�Qz��T	�ڕNX������@���8v�<?4��b��5!�s��"��4h�!��c��/s�y:�
|y�K,�O�G�h1"��MA%|����iq�'��f=���,B2#�J��G5����ρ;�g�c}�Z�'v;���!�c����#켥��l��� ���|�-O�ہ��2Ԓd�R��!TS�m;�1��ga3טX a���H��r�������wWը��y�=Q��k��G9(�>���gTzR���q}����5���x���3�s�XlxVHYEB    cc3b    16b0&��7�ְXu=��AzM'Ŧ��6h�5�QX�}ݢ(,rh����FX��� �	X�L�/ �~'��qe�iئ�;W��(��6.�K/�,�uO�hғfu�>�l͗�kw!�c�����f �r(����n���5�����}$V�`��{�Y��F�Õ�ֺ���N�+�v�ھ�m�G�+�^�:�^�h����3�F��5cr~��A�X����gf�^O.�R�YR����� �7��/�M��oïV���^C�����s�����6%�̚C�j�С�7��@S���⌝�,�Xjt̐�_��{1�S�NWd�>�7�שϳ6!��׃�+wd���w�u�
#A�+��pk(_o���Mۗ�cmP
���j�_n\�?DPL���?�"��t����$zq�����$fK��!�⯾����s�й��r�
��@ap�9ysy�?�8�[i,K�,��ٙSk{�nn�M������� �_w}�B!�u!&*��kvO��g�-
�q��\4$S�V���}�rF�s'fUq
��N���z���0����f�g��!&��9 C_��ܯ�b���.��n�#��jk��dcn_=n��4���!�~�Ӣ�?7�m(��V'b�N����(�3k st�6�g�W�����5���=�)
Tdg�8����"�ad��A�����WD�5����t�N_��"~��,$0ƿu�ò)�#ya'M��B˖��Y�cw�זl&̡hE��%��d�iSM8���ľ)�{n��*fF�L��������.�gv�H�J��U���?H�o �f��{W$�O���'�;@�ǟ��&��}��)�#��H����3۠�9�̑�.1���~/�2o�=LF��B��H�������y�	ڶ��̦zF���X��j��W�=�`H��<�DJ~��!�۔��H؟&�F�?�_!�GHw)�c �q��cw=A�Ց�O���馎���^���q6ݱ/��<l�B��4Կ��h��Τ�8���R2t��-�+p���HLx,5JSZ����W���;�n��1��$N���h$��@����Z�`�g��$'H�<��Tf�½���-2	B�s|B����3b����huή4?h�U��������A=WC?fxg�:���{�@�����.����>b�%��������˒����� �xž�u�m�^�Ou��� G�JTrvk�|�|�z�|� m��@`����ݸ����-��/�\��=�Az;����E���pM�62����RW�-�>����t�?�<8�s`��Y~�G���P{�lv�3q�v�C�8�LzB���+>���rɏ�ߑgv/���ϔ�&t��IuoMx���
�^Yb�#u4�&���m�U쀷�n���rAU^�H��˨��?	�Lh��+t`�����T|*��D��c��6aܗL\�oC�QL���'4�o(�YRx�%����[�a�;+�
&L��q�@Q��1��F(�Rˢ�?��%6�
��� �$K^-�'���R�*gbJ��w���N����6Ƀ@xV�&g#DK��\�2�ur��8��F��B��r��F<z�>�a���7�v�����6RjV�$Ʀ�#����(%Ǥ��А����a����tU��};jm�r��t-:���	��3��
��B�टi��R��a���W�pͣVA��}�����������U����.
�q�i��%VW5��@��V��ҋ�Ԑ�dFM^K���a�a��?%��2��z��l+<k���ݗ@ �v����tcl^Ͷ��i�hٵna��\aٸ�˴ZI3/�j��`p���h�����)��1�9���.{����b�J�4��V������ۊd�Mk�����������2��t/�kO39��$�'��)����X�!�0ǥBU���'���ע{�ð��L-�sZ�:���߬T����o��c�?����?_`<}�T|�yv ����`��5Y�I%"*96�:��o��c8��9���&�z��qEJ'X¼�y���)��J?P��ڬ�/B���pZ�-�0�x�x��5�n��&����
�ljޝbTu:MT�
)<��Bjw�|>c��|�fC�0��dkjKu��A!���wFͅ#�j�ύ7��3�S�K��(�Ŭ��6¡)�^_��w��q�=�Z�����g���ȟ�2�D��Ǵ��[�xI������@�B0�9dD�'Js<����cTL�H�;\_���AF�*��OӜZn���H=�t?�L��C�����w���W�2�9iVk9�d]��ɨ6�����fbcZ�t�%�k\�z����t��J�}l9���	���lE��ߺC�3|���_Z�-��,lIi�u�R����\�E�듣)�޽'w�"���ߺ�@x���.��Yf�J�>����bc\��L�)&2N�M����*��Cκ�$�8�ǉ��Ì%Ӓ���rJ� 7�嘖l����/��=���2�b����C�t��֖�9U���P�Ξ�q<�����D�!E}��렷o�RI��|���#�].�,�vV�D�0�Ck�BU���s�n�R����<�O�T��3"�U��/��ܰTa^b	EDA��ւ�C��"��ՙ��z�j�s�<���=�8%q�O�=�J���vܰ�+�kK��o�?����R�jA�dx�E�g�>_j�0�V�������T�	#b!ʻ�X�I�KsA�t�7zo�2�P�h�d< ��\z)��-H-B�
Аi����(��!�
��}�TR�Ȱei��>-��M�L�ߊ����·Җ5���P:tވD�<ZX7�  ��`�ɝ���*
�X�(,��a���$�hQ�i-�u��c�)�p�*�ܡⰃ~�UD�t�ȭ�}��"%�=�VG�3Y��D�XK�z��o�� 9�Z�&�X�u8�H����.��B�m��߸Y/[�s�μS�x�����_������Aj��3%�ໄ��5������ȏ`��V"�&׿O`e�<�8	�A��_5�J�ż$���0=�1����/�
��dۛj4�#c:(�_��s�LH�m`(
5;ٹʷ�FŜ�z� �y�l����$�h{��q?��6�$��d�����h�GpQ1��[�<���Q�>L���O���j6�I[�kP��Ѯ&�����M6�-��\rIg,���F���������]S�߻���r��?!`d�⺎�.R�>�MYX������ 1�&}�$"��F��05������lI�Ò�%�� o'�
���Z���m�8� ��}�V$� lR��yF�U����H5�����I�g ݦ�~ENi�JQj
�#�6	~g�B�:���ML��,!�hAqZ�0�򥃘i�/(Q���f�@�QʘDp�g��.[�̤��������-�>���#�8�b��Tۣ� ��,�L11�o:��ٸ���[��u��˝�;&��+OaD���Iwi88�>�F8��5e�W��'j%�+��i�f[;3�V���9N�@\_�5@��"��e|*����L%�.}��ƶ�}��g��%�i�3�	o؜6�~sd�q��ZP�1��(��P�Av+�l�t�b�م�j��jE�|�+Fʙ��H��b�~E��T��ԡ�2�G���qRt���jD���4k��Ij�3�*s����a��0R�V+��V��؁�?����S!�X����v4�)%��Z��K�	�z�.�Ũy�W��k�]+&W�=�@��ј��%�0��l��.�A��L���v�gdn�eSyO�>�!Y���vb���$�HF��(sY6�j3�0ǰ\c�Cm��t"9D���d,��FV�`��kË��;�`�gT�|ZAz�;⮳(���=���2�o`��-�珞'�wn۝���x{U�T�m�K�!�h-�*(]�F�͸�� )p����6�sdjpu2�0�fW����{��I�t�bʟ"7E��uS}t�*GZh��h�<i,/i�ު��Xf��æ�憉����������sJj~���1~sN�Q�;ˇ��'��?-v���	ι�~WpJѧ�&�X�]W�q�XnBp��)f��f��#g^�:E!>)�QM�xV�^���-�-9Zd�*���v�<�͌۫��y��̧���@����e�Tk9����Z���Q�Ϭf�6�'���j�Uf�d�����(�!M�/ZkWu�{|d��XD5�bb���Rk�-�=�wn�R����HX����^5�`����(Vh�$x5j�F�lN�~lG�Iь����>�J��R��t��Zb������,��3��8{�77#���>#�I5�?�#$ ��*l�*6�Ig��*���f"��*�r���{�|o�p.�|k�^{n��*��ră�7�mt��8R��\ø��W����v�<!a/$>q�^���ݧ`�~�ֆL'�p5��x�v�#�Yo۶��'�B̰���(�z�����ro/��+�Y�F��D�����
L_"!կ���LY,\�6����[�iu�V�&
����f�cM���ks����),D$��@�:H����A2>���/ǆ��\����h�ЋĎZww֒Ί"m��Eyi�7��<2�TD�e�J�*��6��{��
��)%��Qun�>&n����j���~}�� ԈCv�+�F}�s� ���EE�cqX;���'�p�֖
�gy���v�f�G�m���=�&�R�&uR��D#��T&�c�C�/�h�O�'B����qM��9�E$g�B�UwŎ���+@�>��w�_�k5�Z����.�q+«��;@f ~��% �_�$�a3�5CVE}�c�%�&H/k�(�&;S&D�O�ɥ���gD>���ev%1G����
�E�G>~!�{���Od��B�l;�sH5|D������J��<4q�y�Z��Mӿ�
����ڔ�a��9_��>��^�������hЫ¡/�؃��L{�o�����_���I#T�p%���2pz�X�L�����JPG̬�����`�G��b��3�n|ՙc0����<y^k�3�n�P�_� t Q\V�"=�1��f�KC��KH��(t��'"�p�J؞SL��_F� ��L'�����_m���3 �~��}��>y�IM�Ί�%V��ݴS�(�M���9C](�k"��� �����@���~�Wޏp~�����t��#j�8�(</���n�y���}w�!d7�nh]=_+p���T����܉a��>ߔb�;����̉��^�n��é�70��0���;f��fSs8M��r{F� �i�ɣΆ��6�lF�`�m?��;d�V.�@Z���I�~�J��C-\!�Ĵ����$�ҽ/��	_�a۠�ϸ�~��RX�!(��5�p��'���}9�y	���]B�!^p
�P������� lU�Ug���5"e�UJAu�׸����ƦӘ�z����gU�=�9�2�?�'��K�Ej�vjߟ�T�=�/7^߆Vd�۲������ 8f�7R�O-���
N�m�W+�R�K8�j���1l��] ԅ�B��t2<�z�G�u!���1����k`��%0��x*&�ӌXީ<\[w%��� �ц�zJ�t�bP��ƌ�Eڜ2��G%ڟF�T�;"�zx���Y��VV� �,�