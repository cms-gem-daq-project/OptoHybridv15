XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���pa_�8~/w�aJ�����X�Ht� ��8����L`e��Z_Ps�0���zM��@%�qC��W�%} �������C�/�Ґ(��k�ؙC��J���ڏP���8�SK�1�%]6$ڛ�`��O`q"�I,��\ߑ��ǘ����c��YND$ Z�_�9��^c�������
�Q 1˺k��m���J��o0�G�ݝ*�C��Ro�z�>��.%ب��]�V��t2�j'�Dl������yc�)�$��B(��AeȒ������k�U�zr�[(���+���T�PE9'C��a#�#v~U/��S J�#�w �R��G��m��@&��F��64D7N�ɳUD���~}��N�c��0_���ܴA@�SО9Q!N�ZX[
{)J������o�1�i�'��;�.���k i���9q˪#�R��c��r����޴�=؁�o6�(E��`�P�{R*�\V��8��,���!$���2c����|�|��PKE���Y�  S��#C���b�#��)?>\�� ������!`n������ �曩*����7���j�E���|���~v>�7[�<����<g�'T��횀�6�5�t	u/.��ng�i��i��������}
���ccT��P�=)�9�7�,$�k����d@�e����fvA�X���(ό�XC�mY�k+ 2)mOK@x��ؽUV4�N��՜~��"��Z���1����)P�f�(�淿e�]�=T��$j�Fhl4s*��d���Ϛ�XlxVHYEB    26e0     820-�����Ȥ���h3)�0(�Ʋ^Gr���	F�d���_"��r��?�тl��������!�}�mlt�Z�WG�w�񓉤�j*U�.�GN��bw�^+>�B���+�Q��R6��\�9gr�A�>m>��ԋ�zk�dKD�g��EU��j�j��Kx�ϳ�����hE�m_�Z�ڥ��TR[t��N8��`9U��zby���s�CL|9#@6���^X���ِ(Y����jtrrj2f�O���9#��c�h?�&g�r�"3R�E�쌬�<X�ӄA��b���޿9����<��NS
���f�㪞pX�B�*=*����{�Bnwc�@֧�8N��;���{i���j��a٨��LQD�}i�q����I����E��]����ܾ��_0'=�K,��Ф��/����[l:3��R��3�����b�0;��{������s�,@�� �;J��rD���'bS�@�T�?޷�/k�I���.GE%��������O�v$R��P�� �2�&�2Z�d�@S)R*��cm��G��i��ù�QM��y�_�qǋ���R����kUU����,V�V��	[����*�V�0(9�^���v�S�|��Jğ뗝2_���l�kG����q9$Mxek�C�;
\m��C4��Q�����yh�F}�f��)���\�`��XY���3Xo�h�2֯s�yN{ �:���������ێ�1Ygq�%�F<�ϡp~��̟�q����?m�]�h�Es��免���>����Cv��ᙺ����8�d�5.j�Rֲ�5�=��'�	.��.�ޏ�	-����c=��j.<䯔��U�F���K� �֒ ���z/B���Y��v�n��]$���ۃ����a*_>���,ܶ����^��d:S4�M�٣��Sxܶ�皜N�;�.	���K�1B�H���[:­�r.칰aE�����P�ST��n�B�_��y�z�d����Q\M�י��&1�ó0����
У��a�F��,nkt-H��Ĩ�<���sS�%��>��le8��FeB�Q�In'�&{��_�T(Q7V��(�l���/�N������+�s'Rg��y_�F.'$ ���c��h#]��yj;�����o�۴W��D�~�#4=�;w:� as�t�����֢���6�i��+U�/��8@ψ;�8��K��249Hf��LH8z�.c犲1̓���nۋ�e���qM]	��$����%!u�I�m�"�M��R���%)�ވ|�h$�,�;_aQ���]��ӑ�AJ�nu�Pl�u�|�f�7��톗1�p��=60�����$��[!��d�ʸH3f�?�H�	�:KM���0��S����jy��7�u��ꯄ�PjyKo������z\l���&���%��x(���W��/>ˈ�	�x�����-t��&N�7)�xߦ\���MR�h���v�X��:���F�`d�Ołi�+�ɬ]�+*�ԉ8D�h�hmۥ��;�u�29)Fd����Y�ү`!f+�	�"e"`�4�үS(2Jb��tP)G.�p���p	�MO���6A������V�ƛ��v�|�:��,W����� �v�U��j�5� <��r�`*$3B\�m�9��6��a�o�M U�+��(���J��p�G�o%�e�:�f%����O��Lb������sGRK���e
�w텠�k�����NW�=fu����8�X�V:�3*L��1/QR4���w}���Y�ƞ��0����Ο�)��7���ڨ"�YBx���P�1G��ф�vG2j6ҌC�\�c���< ��+hI��[LԾ���&�e��/��m5��j�㊄)��+�A��� ��#z���Zy)ǋ����`�Vm��sK��P6���A��9��4ݹ�*`a��	��E���7}TBaj	>;G��ո4�tF��SQh���~�h��la��t�_��sG�2����KH|�A�	��kz@DЇ�=�O�l	tzԣ�Y|�ą�L�[{�MZ+��s5ѯd�,"�j��