XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�sV,ט���_�h@G���71D�D�d��{���ʹk���� �p�N����!��U�9��Y	���&P- 5���J#~���> 峏�i:��r��,�a�mK��o�����_DEd�YA�}�Gv����9�Qh�V�xq;Nh'�)��^��K�|��d�O�����DZ�YO�"/V�0������!:�[q����n�Kw6ڮq>��w��	U�AzA)�����4�,:��"���%��2>�����h���b���W���%R[���и�j�|}I
��	�Ѯ_x�oq�7J�f%t��ml�L%�b�C����&���=�����^s���o�Ǝ�	<�%�s{����xbԤ�xй�eu����d��F"Ly��l�03/���L��C��(�"���)^y/k�wLO�YlΪ~�}���;���O3����ڤ�9���������M����$ i݂s������8��<��A�RQ��X��T��T�))�'�nKS�zZR�2Q�N׌�L���M�c,	* ��]v�i�Ô���A*k]�)���R	=��!(m�(�C[������,�����jNK/cg�^�O� 뫂k�e.B��Lƙg��zY��.�ۉ{�r�y;��T��r�S`X�,xM��%#9v�p����m������D�Q�B��Z�����Zbڣ��ɯ�j�3h�\oKv�-ɫ���	�
�ʺzKx��k���c+��#�mP0f촅�kUXlxVHYEB    1047     4a0�eX�a��w(�4���f뙚��fэ3��0]2dg|�c��s����o�B]t:8jk�*!����"s�m+���Q�3Y� -��GlOV�	�W�9E��� ^���	X)oO�p����p(:W�I��'�h�5H��yQ�EZ�'��ľ��m �.hJK,Cj�3n��4��oQ��5
�������hR����;�e�BrbQ����no�>����L�F�|���|J9_[���ɲIS��D^�Y�V��#l��H�UJm
�?{�`���@.�N#߹�K<©�{~��bͷ/U+�D�]��ȋ�dυM�lgH��׆J�5���ʞ�U���a4t�(�;/�9��E'U�6jF�y6$�����C(�����=ʜ5�#����q�{�4�?w�B	��$�Z5�"x*$�^�����L���m��� '�ts��y��2���߻p���`2N��Peem�{xR��t��c`�M:^�/ߺN�M=L�F�!��Ѡ𥝨��em���P������{d|�Μ�J�E��ugk&�S�HO�ŰU�U�,ǉ�'�{v�뤧�1yg-�3��=^���F�m����_�-U�	JH�U�X{@c�΢L��s�ߟ�$jv��(� x�,(�F�/P�6��Q_Y��{�̺j=����V�-Tj p5�������4l�����t�Fl��h8L?�'ҟ����}�.�TuU��$fX����:z������.#���b��/�'�.�3��'�E��΃6�+!2@��(q���-5�j���X�t��:#(���O�	��;�c��}cuh��
�1U�;K+ФJ,rsq��6Y������Q�U:���c���� |1��ГW����趟�-����m�IG5(�ņ��MP�sk�p�Fh&�ҭ�a�t��@��r�$�Ⳙ?w��"M�tV��!5x���/�2�=Sl�<���Cd	!�j��#�W�������=�N9k�-���&�(�j�)�cF�V4@�9�Y�&J����
�EؓȭJ[
{��ǁ9:;�4*��	 d9��4`J�%��w??����YX_\����Ei�h�AXjM��Ōv��g�涁��$#z���&��CaLDm�� �H������0W�z���q m��-X/>�O