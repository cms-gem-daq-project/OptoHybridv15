XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����5����2dr������5��� 8����Onx�"!� ��Z�:��x@��NG��"���T&}�9���ʞ�1����������(i���g�D�7,#�D���#�sħ��*�Y>"�e�e��q�P등�`�۫`&������j�H���:�A;2��&��Y����4�7&&��<b�+g�d�:3U�^0�Ψ+XO%KE�ON��C~�[F*�	��g'r��~6�D4M�F5!Lw���'*��aR- sq��JL�_��S�L�|(�f��@B�'�|��2ϲUr�?�%֨l�`�e�-"��hxD�z9�V��$��� ���`� ��Ԙ�g҅��9f돩�/	�b�̰��6(�K�s����z" �Z�0� �>�S����1*f"���͛�}�5����#+b��L
Q�rz�r��5�; g�+��$*-��5�/�m������{���N?u>J�_����kM�4�a�Kd��
@�K�d(e&�ٿf�C� �C��<S�����mn�����p�6t뚌���D�O .����?u�����a����h���ExkOW:��^,���U8���پ4<�0�N�B(M��y��b���l�A����|a�L��*zU]𦔐�~�u�`�y�>J.m����U��6Ƙ�KB:r�t����[�;����V }��ǁM�֟��4j63�A�� LW\Dx_>�S�_��?0A��*P�G�w�e�?A��*8��pXlxVHYEB    1046     4a0�Z���
�ۄ���8+�D<q�y��^���*�J@�i�yăՑ��ˆ����WSZ�C��D��N��V�5�J�l��OHt�D���rq[U�0���`�k�m̅E��.��Y$���/�1i�0���\)(-�^\�f���yO�8�'�V�o��(��:�̮�:Ry������z�P�u<F�����7�����f[�5�Fx�SIG���7��y6�}4�|L+�%
����*,�П�s�	�YV�>��ز+������;NxcM8,��D>j�V�>2�rE����W��/������Q��jF��ɲ�t9�?1��_��@4a���%t�S�FS(�K�AuH�7�A�|A���L��&��~_ེ���hl��?IH�I���j6� �������:w=B��_Ы�>�n'n�=���h���L��S���Ws��]x��a�7�25Y�
�b���XS�+l��d&�I�v�6W6l�� �C����-�i�O�@~�I����T���0���,�96�I�	�h%08��k�'�.�ۊK� �V���XH�	��9��1^R�#�7ޕ�����8�f���q�=$4?\���g���Z�lvf@#6��.I�Dp$X[o��} V����s�^�*5a����ZԺߺ�P�R�9Ӡ��h<Aꔍ�P}��������ŽC|	��/��I6�k����I��ӻE�Kx��Q����ᣋB� �S�l����r�A�R�id�F�|�t�b����'��7�z�B���y�/I���	FD^���F�5F�F_WQBV��D~����lQO�9۳��L&��Z�Q����7�� ;�u�5�4��c�S�5�p��'WOIzX �Y��ac��.VG�=���o�L�
e5��	��b!�����ќ���M�f9X_"��%����'�ŶE8�e���H܋y�1!���d���ݹ\MG�-X|*j�)���b؟`����z��=a�v.�N�������R1?�_�ocᢨyV�퇑\�/�A�@� Qߖ�Sy|=�"���aP1L&Z�_T����B�e�.R�Ś+wbJ?gFs73B�܉����#��=�l��E<�X�<e�q�d_��t�2�5撧����6�ݳqCɠgS���L&�ļ�
�����,�,�V滖��AJ� e����٥A�P�x�k�o�'