XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#ׂ�e/hm�cO0�/E�7�2XV�����k��\��^]�_��X�Q��	�O��ۤ�s�{�ov�E-e�$�k��6�^_�2�MC(3-:c�]��&
�Cþx yM.a�����Ŕ�ݱ�tVW�X��zf�W�zl�������4�����#�����S%��*Т�����%74�8R-�d���w'�)�F��Vլ�K�������Ǜ�SUYA�����Q����eA�]%�O��WXv���.},��%�Ɣv'�S۽e�Y�M<�?�NS���=o����1�5БSB��`qi��Q��M�y�&�
fQ�<o5���,ӱ�@r3-:�h��E���j4�Z�(4�U->���H�A}��mq{���*-C�5��<��
���'�"ojh��Qד�TpU/� w0j�̳�o5�S��T�Y���43%m�����'Y'U�	hqHz����6���B��|�u����kѓ"U ��d�쁢L4��=�]������3�I5͡��c�e+Y��x	�L�cd�X��/�vwjv�|�]cܧ6�SzЌfğ�+�y��D�<A��J�����ͷ����k�͕����)naf�	Ì�(��ƿ^x�i5������xH���Z'��)�9��Y���n|&�8�ӫ��ъ����4�+��C���	���j�ݙ���,��uD w!�zM��#p���ES�Ճ�K�C�r�C�FP�.>�=:w�<4�([0<�����Tm�}XlxVHYEB    3c90     900��*f��@_i:z��z���t�M�\wKS���Xg��Y1�5c�Mgy^�8a�AZ�X����*�ks>D3�>���ېN��c!M8��
��6�)�7�;�ΥI�����Q%��]�Y�HP�N��~`�ս��߿��8Urgi^g��fk�F�O��03��2 +�u�ް��YKj�1
p���~P[��H�Gw^O����)U��ʢ5-���p9��7�:RH��2h�9��!:�]���A�W���qC�6����t�����F(���G�n��6��J%�Ⱥ�-�V�U�t<�q5kX"}��#hW�x?eN�гF*���8:�qvau�OF��<��N�0�Z�0�=�G��˻��s�;ғ��~�`��^m5��f@UC��(�O�m"yn������\�W�+��R���Q$B �����ft��L�d�X. oD�LuD{�p���I�a�of�E��W�+����D��?	�Nd�aWj��-��a�zJ�Z�&r���ָx�v���մ��3�T�>���NT$��b�6��(�O�;��n��+;IN`S�~�O[^;�KFLi�([�����i�T���<�Q�2���3��x=��9b=0ZM�NkQ�MjGi�B���4��a�q�R1�ɲ;�,��ϴq�~Y�`%�dC�H?Gc,��Q�}&i��s�RD��ҝQȜ���7�O_��RәZ��d�=�ҍeq$n���F�����e-9�&w}��@נ�f�]B��ҋ~�U%1�>� ޶�un,fge�zŐi��m�͑��Em<!���F���;����7S��7+ A}��L���4J��2�ecl�9�^�2�b�l�L��+V������i�����,��P��W�]�@���C��~����б���� �{�HQoL�1C*���?���͆��Q����J���Kn����|_��&^f���Eݕ:$n�9�k:��g���O8��^�*�~Z����0V�J�kq3h���]Ei� �)�A��#�_�^ H���m �;'�U�
�|_��kH�y�cR��^js��6�� sa����F�e�j�.���N���z�7�C!{�R��"��3����;��<c;�T6m�Mx��w����kՁ	a|;�1l�6�B�C#!���с iAlw�3�@'A7V�va�;v����F܄�o<�A� %��U߾���,��A���cw/T��/]Q��u�-ɪCQ���8LA[���Ѵ~��T�@KgE4q�V�T}��3'dR�ܮ��L���=!T7����G��� \�N�P�.�r]Q7Z����$�6\����1>,���M���@�v]��%�;a�@v�U�w���Ο*��E�z3�0e.=�E]5�p";e�YU��gk�O�"K ��.���%r}�Ism�'����ת�C�����f7�bWasS����� �CYT�T���;���4O���A~�g�>󗣫�+G�X��=��[^��P�~p�ѷ��9������v��6���ꌓP�}�A�Mz�L<�#���˚Gr֟5�!Mu�t�PQ���P���IiB�.h��O �+����1n)s�\j����ny�oY�y%�q��Loh�V❽β�fN���O��x9�W ��F�@��7?�zg��Ͱ�SRP��N����ڄ̙����5�u�̤�FX����	�!*!p%��2��c����¶!�>���30MA�P¢f��%�P��dm���KMcy�fr�^�]a�j���ܭ)��Z{�M�E�O�vw�c�H^�К��/p:1�s��y��Hhp~�g2�9�� ]|K2����d�W�ϖɩ��C$�`V{�y�5CY�D7CP������ ������H4��f�,H��������Ӱv]Z��g�����@�Z}$�ab1������뚐"����;�J�hKH$��G$ep��-�r[f2�3�$a�����O�-����K���z��ۆ����Lԍ�7�pA��]��#0�8u�"��Q��cߵKl�i�&iG�Y469�zFf	���e/����0ǲz[���4�@U^���ճE`Җ/�(--�vB�3��H�?�%0mp��g�>8��h$MXLF��y�I< :Jm� ��=V-��;ϼ&��j⹪��7�2Y��}+��g����w� ߓK����6<���V�=e��prXc�ڻ���hoh��s��C�Җ5���^�������Y�(Z��Ϯ