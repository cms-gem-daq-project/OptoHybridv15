XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�0�f҃=RD�ÒBR�+����k�+��+�H2�l����e��`�\>D�����i�[0�=�-�mI^��	Y���Ѣ��M�&^���a��U%gP��"��9v>b�Ml"��

X��sg�PQ����X����Ǧ����2eu�}�0�V�KԲ�i���4����{�c��˻�㚟��V�l���t�T��P\�-��w��/�>��Ƒ}�w��H)Հ������hEw�˶ț��lb</Jq>�{�s	�������Ǹ������so��<�"�ϐ��glڦ��[�{m�TCLGI�@�g=w���Έ%x��蕕��H"�Hwr�)��1�fe(�Z�����z�,6���d��.��+��&ӚV��S����܋�^����{si�����S�k�)���΀�g�sՇ�Q^�a.��_��`_H�:��ǻ�Y���"���2!�r�MԱhZ�W�tT���Au-:�l]5�~η�h�PA�Å��ˤ���S9�K��U?rʬK�]��7#(�+�a`3Sfwͮ=�MU�JZo��/� ����u��k��q��fE!O�i��ؙ��suu�v�64�G8����o��)S em��u���B�Ic�/��lԩ��-�a�=����j�\6�;�����C�/Zc!�E^$7�E��ywcvˢ.��!�@PV�"X3UJ��7��S��==\8=��k��zX`��="֡��:xK+/|QC���Q����bu&wc`����cz�XlxVHYEB    5ff4    1040 S3+��F�k���x�=N�qc��)�RRUe����9�P�6n:�6�1*�XF9�A�Ґ@FK�q0�UFYvW0�辙y��1mv9V��"��{��h�sX������I0�C��jLcy��Nm:�pB�Q��?�:�e�R;Tf���Bӎ=�l`OD��8m�f��u�Z筢j��X$�<�8�ߣ �"1s8��[Mؿ�BZ�{�	Y���í$W�O��Pj��o�B�|��ɶu"ny<.ʅ�P5D��:�y< ��2Wt����YߺUt����څ�dmUQ("|s��*�L»
�L>�ɲF�5^ɦGI8�ш#�ҙG3n�Ǣ�n{Bcc@=D|����f�s-��k���L�^BB|�z<o�_�G�0���`���|��\�Z��^�4l�v��>�p�8�'����w�Ӎ�eJ��
-w)�́=	mJ�+��X~�̨\ND/*e.����1��U>ΪќD"��7'st�j�m�O`��|�,�= U���`ߊw��9�ē[r"�r�ʰ����|e�����1�_Zނ�R��ź�Q%R5h�l�Fb*�5?���lVWW�U��th�����vY%S�T�p�Zq�`{�"<��6N�1P�1 ��!���ҟ�F�������ʄė<��ۉ-�z�c8>�N��Lv@��&P'_�ZV\���ò��+Ia�y��5|�1HUQ�p����֛�C�;6ABF�]�m�Z}�tSJ|�Z	cQL��4XL�Y�vVT+!��8#I�v̯���������#DUe�j3�]���<�C�%lO0��,�ƹ��(l�tDE�m�6�Puk2Ǫ�}��u7>��+�u4ޢ��(�yκrtr�:}9cg3�/&��İX.�7x�>T�׊��ι��;p�:/L�]MB7�v�+l��ۘ���ۈ�����4O��,xjB�e'/�Юv�Դ���D�A��{�*
VQ\�n�K��@:�:����wH�X�	�����OO��|Z���H9ss�_/�Y*m�ARD�CZԠ�I+��L�*��4w�8?7c��'����AKR!_!Q��W��'m�948���8�(S���I�\2R���&��ݔ²]
��^�"��ܠ�x
���s��Aݚa��7�H_OM�q���Z!��qɪ�KIZ�C,����6�2��"Tj׺���s�v�i*C�7{�>���#��Ǌ������ccŸ:�B���*��%��Kd��p��Vo��M����!F��\uB�ɂ[����M'�}�ᒲD�blI��U���0�|�.q�ɚ�-�6�p��!o'�z�Lu��`�{I�#\�l�(�}\�\�p�6��a��N���.�S�d�OZv%f؂�gA��MS�W��(s��$�%"����φ%D`_M�s�y�2�u�y���HB�����a��K���~Kh����#���[��'P!?�Tܴ�ƇP7[��������iii��G�T쥼���G�7|�Ġ�:�{c?T��H�R�P���e�tK]:NZqS/���xЌ��.}��Wk���Y��/V䡅��!2!�V�00�I���^\ڟ�&ܓI��fC�.����q֊�.zB�K�.�d7"�j��b��[jƲ���k�)7;�5O�E����߁	#(�:s2_[e_���P�}�}H�1���=�g��%��&��v��ܹ�=p�����I۱�i<���_y|�h���j �3�q�!W�د�T9QG���`��/�S�b�D�p���}�����Vo�;�VM`���F�>''���G�3��s�6�5�A�i��S<S5�k��8&��p3/#���՛
g��P:��y᭍��a��]�ړ�[�?3n�}�� r�	tW�|u(�m����Goj�Y��r��^�F��S�\�٨,��j)�<}u%=c�:���C�" �f⇣���4��w��E�W�v���$i�miC���>�dHB�`��+�J}S��L����,M�*�f!����@����h�/"��qk�b-V�3��<օ�<R�l�?V�ןe%C79�p�,�TS�m��S\�׸�u=�����}k�9�x��L�Ւx�e!�3���S@&����ƪѦ\��z)R�6m(�b�W�},XSYUr6W'�z�t�WV{LF��CI��x����b��*U��x<�v�3��Sn�\���Lq�1Z��lu,,4�U�K����@ʼ���>x�Ĺ�L���+��gi��ch��U.O>}�o��lO�%^�5ߎ`)qe}�����~׷��Y�ї9�OU�>�]� �k��k*+��n��Br<"���:�?FjO'��7i�U��!�T���PPW<'ˬ���DO�WF�Yr���vO��o��Cc�>;S�����4�k���C�g���t�=���>��ۘn���W��H����,��8S��!��|��I3z:���@����#:x�����֪��D�0O�4��#)�NI����`�Ă���S-e��_��v
,ՈK�7LT>�	��z-*�m���b���.�>�^�D?�_W�ݒ�Z%�*G$��O�6�5����	�[gJ����Pԭ �&�����,z�'_�Lṉ��Y�$�~�1U���9�g�95")E'ۏ+={1�Z��#��~� ���(LaM+H�.��2 9~��:�%b��ft�BU�)��(��I4�絞8U?�X�&~��<&�8�-�t �E� �x�'�*�����S8���&�*��2���,��`�$�?��>v��+���߀ ��wF}G��L'!U|�U'�{ʠ��H�#� P�HYd�#�^ '�vm��� �F2'�qg6Hg;`ve:X��P���v椟=��3��� bu��!$A����5ײ�3��*�R_�]��-�UӉ�����Sp`��%wRN�L��̊��!Ǯ��,B�e�ա���O7��l+�e���7U��[ڤ6��b�fG����
��g;x+��΀h�����BH%�8l/�����t���Uߕ��n�\�f#FR;��D��d�C��#a�|�3z
�7�Z��O1�?�,9Bcbn̼�ث�4q(���Y�(L���ha�9yֺ��Zd�����1}�PǠ���	zy�E��*�a2	��O�.C&M&�C�<�����phư{�R�	��Cߓ������ m������U�Dl	&nU�X>��9J+h�\x_WJ��=�%��_��.��l%m\�b=��Z%�z=��	�!���{O��G�|�������ww$��H�҄`���$�Smԯ*�� p�p�}�e�J>��H;7<z��+y &R����T��g�-ٲ��[U^}��%W����D~ι�If7�b=j��T�+�Cs�������ut(��N��<<HwL��*��s�um�n�&�!����6�G�Idi&Pr�t��2�������� ��M؋#}2W���m:.Fv@��� `c�n���JN�)��q� 6�^q`'��Yo�/qBcjT=��"u���d],!48�>\�J�:�G�Н,ogUioUF��ii:�
��T鯯)c$93���w��0�ڽA]���m���J�ˍ�c���p�Ϲ��}NO�R<N�a���Ò}Um拃I
�C$���s R�kv��"N��Vsp��
l�p�#�tQB��F�s���n�;�a�`)\,q����k�<	�d�I�ҽ�LI��'ST9���C�����}�����.���c0j��G��?��j^]��-0�E[��Y�k���� ι�Π��n��fR� ��Q��d�vvX-��4�F9��p���/t�N<�,{�5+t�dχ�eP�_a}5��W���<+w��\�����}j8A��y{��ф��Qϫ��a.F�����?�͕�E˳?]G�}���i���2ǟ�!qd�OH .�ڹhc������!ϝup��������!R&~�bZc*v-���x�G5�[sA��kEV*�e�F�\���lz}�"*c��t#>3���r�`ɩ��:h�l�k�΋g�������{��2�M�DH��q_�.��(Y�����#tK�|�Mr6�[o��6�o��S