XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AX�?��^�y�tq3�u�E�[�W`�&�?�'ڤ�D������UV?L`�>ݼ?P�dk�A�'��ю��m����&�l�� �<20���mL:t� 1����Q`]=����f7N/:���U��o�s�l�UV�^z�L�;����K��x�;�$=P}���d�5��(%E��ႚy��(��0׃c�;��߈����r}b)1L�q4�x
���q�3B�g�C�:�y�[n�j]`�F�Zz?�l���h��h�3>��
�Io�4ܱ�nVtK&��X���a�育���ƾ6��.�4N"w�]�>�jb(XS�S�������q~�z$�D?[���uS�Br2��V[{y�
��:�Gf�M�Jos`�mL��5��FI*
7��@
�U���F15�S`���ͧ�����`�L�?)Y1WIx锲�/jґ�*T��bߛ�� �MK�Ҕk���xS,�T�8��H���_���.�/�8r�r���8K��zv�k����k���-d�:�n��C'u��n�!̣-�b"��$�R2���9��:Q�w�k���KN�V
�7���*�f�g�m��p&���5������o���U�����V�LP��ɠA��y��1n��f\t�yŢ�:��b�L\�|�y��*-OaI��d� Q�����T�E��1��L�d@K�@���[��"��C����Ȁ�μz��`ISf�:��;�c��Js���R��f���\�e&��M��k1�B�u���XlxVHYEB    fa00    1960��,it����QW5�=^�W���79��j�K�Ӆ��k=�z��N������On8��U��(�E�b���#w�0�I��=�l�¬S��0V��b)���e3�0�n�L�Q5=���(e����O���)�PB#��d�(���u#V99�{9i�o&X����������h5��"x:%s�bm�)���ө|�?��cٳ�{����\/�޸���hk���g�"?y�u��B��d3�J�e�+�EEg�'��d�肦��J3I��&����{�U�t\ʸ���*;��Z�ː	w�1�����_z���$7�+MK		�{�a��l�cu����:�<�����f雙#I1����ϕ�����,��fQ����n� ?H3`pq�HGo��d'���;(��z���e?�<-��x�D�3���;V���˰$BM_���|^2��i�Y��Yf���.�����&ZC"�$-�3�s��2�X\	7;�7��U�H6^" ����j����{����S 5�Yn_j E�dn��Ӏ���J���*���'��(�R�pXM���N!�A�/�&�i�p�®`�i>��W���τWA�h,�m���;�܁O����f}j��hh��Kzh7y^$<_$`��52�W�	�;��i}���`)�c}ΕHc���g@�j쾕ݘ�Qėжrք�I!��첚0��,�㸴�U�7y.��@��FOh��o����N/�navN�v~.�^���(A�5RR׉�M;�Q� �P(�v���u9��svp��8Wf���S�'<fd��σi�N��Vg���:��S�Q'ucL����eH�6C�)�9)A|�}�:�L����/Q�n-��	k��R4���1B %��r,��.{9�&;��@iQ��B�C�u
�i�|O����Q�4(P�� �U\����|�5G��QW���Rf��o�=�K(�T�o�8Q�J.���Y��&M�:^XYc��x����m��m��=��/�.d�� �)^#.V4]�RD���h�0_��쑤U޳H�����2xu<�m�oݪ��|�z��\�wp���u��Y��闢p�u�ǚ �ZF9�Jk�̈́ͺY����W4��S�Z4(�z]�)|�� ����,BIa�Y����g�Qf���bJm;.rv�ȅ�Kϱ�r2��Y�FA
�tXɆ(��������L�6g�Q�~gc���^�ā�RP�^�C𗗿[t��α��ǡ8�eq�rs�ݱ��tw�S��譥�r+��$vX.�l �����}����5栃���;����
�.�nɐ��Ϣ~6�Rwsd�j%���PU۽�<�,�{�n��H*�Ū�m�ܼ��?�+�,9[<b���Έ����CH����ʋ��N�Ӓ��r�v�ɒ��E�D�|��[d@�`N@*Ǯ����a�U�"i,��ݢP����u�%`�t��.>;;���F_��r�Hm*��)6����ϣi�����;eA�h�_e2�o�3�����A�_��/������7z���sU���P���Y����9��|�J�J�#��y�_�8��4��ك�օb��dȘ<�����X^z�Xtه��P��QlDc�$��p&y� �M5�Jsb�� cfRc�!����r�Ŏm��]�鿲�]ʤ�����G��4)�����g?���[M�����մB�c�+��M��Uv�崓[̒���?1���=\�~��C
sS��ͪ�:�H1�eX�c��,&�$� ����%��S��#��a��7�<@�=5���s2�>1EJ���_�J�!s��c� ��Qg�[ ����0���k�	���ܡ�ߢ�+-xJ��Dju���}	��v�U�r%$������W���7S��T�e"D�G�&/T;ߙ��>��rҨ�Um8��2� �_?s��*�ٽ�/:���Y-W��Z��&�g'Vr��=-����8�P���5� u�V��^r�c�����N�O@+0}���oB
o���<q霖X�{GWZ<�"u"���[~5���;Gp7������8�6U��K-����z�|�2�5,�S��0R�q�_�{�M����M[�:�����\�Ef-�V�-�lR	�m�G�c��[辟�%���V�_����b]tI�:�]͈
2�a��4��7�P?�˕�o��;���-=�i��4�vʵ�3 �ڗ��z��Z�rNI![?t�L��j�՝k�@��)�T0�� H�T*Lv�m8�QPr� �ޚP)Hd���=Y"�%7{!��^�GR���B����%�w���z�5~p:)�t�U�|��39�я>f�=_�X�xB;T�7Wq-�r���	ɻ������{����k$�Yu/�.b!aR�_hw'�W�g��7ݪ-�t����G2n��ܜ�q$<��py�j�#��1ZS�frJm0=ZN��>߷FlC���d�
f�۶��G��I�����	���eT��]E�!�L�IڲD�pht�gh��SK`�y*E�s��}�{�����|�Ш��W�z�b'G�F�\D5,M\�;�5�~�ʈB����S���7����(���׽�6q����ָ�Z��	�D-���ʠA�aSV2��I�n�{<7BE�w��Zd�'$0�Y ���Qy�V�����/�tE�O���׋�8+-�rX�,�,Z~$�~����7'ҭ��	?H//�lz����u���ը�uk@譙[��I��F�� 98���F��\}N@A
���֌�f���͈��71���]z �D��0��?��p�����#`���|��aW?i�e��8A��כ���Ft�]>J�e�	4�-B��w���G�X�Y�'�g;&��L��l�%[2�� S�)R���7��J������1q.A��9�GOH�1(���~x����S;�w��,,X��M�#���7��Sܛ+8p��ࡷ�,5='�Y������3�ن����9H��yٺYsO�g�u��F�ѐi�C�l��M��x�G���B)EO�l���n�o�������"0���Ǯ�[�<���qu�Ś'�2N����+�~�hӲ��d!��q��z���A���f�G���I��n�Q,_-Wf"
mc��sr�1e:���� )��UJE�!kYN��/5uY����ot��&G��uu�U����Z��٬;���,g�rO%�x�FT����'5;mg�4�gɅw�ǐρ��iC���5E)�Te[��9p�ط�� l��.+�#!�r��A�p*VӬ?�SE�X,F��Yg��tg�a�5���IgM��8ߦ��H��O��Ir#�|����bI!��`��إ�����e�96��m�a���HD%	 ���'*��v��� ��k�mV��U�	�ȃ������-~��*��ȋh�fM���5������U������4ϗp��^��9e��+`_���]�����J����}�zP݊~k��6�Nc�8W����TxT�TE�F8FB�u��S�%8p�Q?,�S8]�1Q�Zs�	Vw��,�vjf�[z�\Z�eO��0)3�a�Ա*˿�F܈R��hV��,6ۢ����?�5�2�_�='��d����� v<	b�,t��PRX��+��n�q"N"Į���� J8�a�DT�K�x�*�Ҥ;#�yW^A�=z���R�������}Kz�#wŬK�ޞs_�&Ʋp����`1-ī@�'Vvդ��L��Y�5����d�'Gq���3��N�c�˭��VV�P�wt���A�;�k�	n��R�*���=�wm�;��hK�l��&�>�*W�E�Hu�*S3���P�:�0�w�u�6r~o��CUж�֯�
��%��8�y�)�D��1�t�	�{�����g�Ew+zE�ȳ��� �m%���P�]��l����ఆ���,��?�RY��l�M�5�J^��NA�7 ��\��cVU6�
IB.��ʿU>�#�˸��3uqq��� ���1��*������n0��%�#zǴ+�ų-�4�YF�l�]+���i�50ʲ�F�vA����}�pi����䝦�j�g�PI����S�y6�<��|�Pp����(���&��d�/`ڮ�����.k��+�qrHo�Y9c�~��1�~�}R�����<��c_?�D��ϔ��������_Cd�ӝN�xm��t��S�nQMP�n�g��;9o���:��-�1���R��[�0Yl]�B��Y�w��׀ּ�9�Ŏ1�:���=g~����o#�@�H9"�|n%-�N�?�����a�+��]����[�l�ԗ�����Vr��\�ňieB��%�݅t�OI��;f믍�!�����ڡj� ��҂<V����	#i�b�0z��7ٗ
n���} ��'�@ik�{~��~��jY�g�o���r�LE�ˏXb�j@�S&�&��%cY�Cֹ�#����a��t�Emz�K"�5wL��H�,	�8��<Og@6��;����T�i��ٯD�B���\�� jb��F�=.�}d^c�Aض�a߀�Y�ŏ��֭H_�m�����D	�,��X�r	���-$�𩞴H����Inr�tkĊ~m��Ֆ�Q�w�����a���=_��ʑޝ�qp��G�V�(Xe8�k�uH17aT�	�Y�#�\�� &B����xu�zt���Ǹ=�!��'>�j���9rtc��m��/�����Ic0{�7лё�iC�M�	�Q��"c���KRX0�aZ�Lx��z�ɼp�,��#qB�V�`$~\5�U�����l�RR�wZq'�V�/�����f��nH?���FKj/��6��6䵵j`��C+�*[��Es��GuIt��%��ue-,�8�m|IX�aQ�W��>��J��FRQ�{L�~��Si=*i(����w�	|��Ȧ㴕ĝG|������½�������F.㠪un�y��Dp��U����Y�m��i����@��M�XO�����)�ы�X�:�k��ϯ�×�xwFnp5k��@6�̄ϓ��Q�������B�])���NzA�k�d����U+��˵�#�?����A�L?M��{�^a��C�C�b�	�~ HLG��^dSJ{�cK�M�1C7/�ڡ�%�p�HI%O~�������-�:�7���&�Yۖ[X2����~�C����,g�HuX��/ӯET��I�D�|G�o��m�*�"Q�7�����{�!)�	��ͯ�8��;�r@��F^C�*����H�[��K�)����~�����X"�����<́�n��Ȯܖ�{�ol1�c��v#�e�B�C/���P�nܬ= �������@Ѣ>�u�dઈ�%=.sW�|j��|�H��(�ȍ�!����.z�7���k��h�3� �Bv���	S��4N�D�A�5������Jfr�8bw�x�V���׸�<-~~nͫt!DOF}_��ɍ�t�%"�l"EG�X�k����
>�؜(PT�����E2�����T37�.X�m��"t1�$3��B�c[����C��)z?Y7ͷ.~A�~�9��;!�k�����Z�ڕ�:���8yEY�(�.x(@��$�ca��a�y�m�%*'�w)�C����p�����=J�����Z%f�v\�_%������V���P8���q��#)Q�m�s��M)-��J�����o�/RgUKiG.��L��N���_C��zv��e��ދӵ�=T��{�P.$�	� ���o�X�Ғ�,�#	7�#�bYG܉�A0:�qw����5����;�������H����R����ɘ��0�Z	���fn�eb�b�+x��rI���P�&�o�C9�JP|ؒ� A
���AV�-P+ą��ܯ^vc��Ծ�(��w	>P#-��u��q����V���d5�H�S�i�(w �PՈ	��r��4x�9+�S#���Q������,���W��p����_���Ȉ#{y,�'Pp:OSM� 6kFY�xDf_��!��
�ܝה|��_ H�c�6_c��f�<+���s����K|
x�1�{�e�2pkGh�����	oM�d��V�?L}ߡgHE0��\ȟ�1H7�[�$��r?D�bڌ��9'l� �j��C㗜�ۊh� �@;�H���V��FX��G)�^�w�{`|34����2��um�'�Q2}'��}u���A� �"J6������W�4\��s"	��&�Gd�5ԃK���6-�P���$s���-7��rNl�A�֬E�W_�ѴqH�K5sv��f
/0+�g�7���\/����G?u[S]�b+�W�U��:�Vҹ�B�ȭJf�gq�P ��8q��˷��8h~nA�z��ӝ #XlxVHYEB    fa00    15b0e\T��_��Ed���;y��T��.b\t�y���9IEw:�}��ID#��<͗��`������Y��_�;R��q�P�!Xfu�����Z[��Ɩ���Oe"�m�0 �k䤺:?\�4�����#N}z"_�/���й�F>��&�Fc(���rf�7�w����0����ZLs��L��Ȋ|�ʮO7��S�\�O#�G8����i}3{�È˖[�m(�Sl-�#[Âlb{9��(-MH�.3ʔ�᪰�յ�[�Hn�VM�5}-EA�=L�����v���Ж󇡘2��َ];b����nF$��޶��z'a���=/���R�������VM5U�P�Q��f?��t�u[�37΋���ūP��_�w�-	b�n��m�TUk�w��d�m&����=a,� Y.�I�m�����&�1p�qj���n��&���`�� ����j������mVz�e��߻p�Ew[�<�z���s��w��qB3��E���H����$m[�'�Qr0�4F���U[_�t[{��u��d(�j�g�%f�_�+� �~�\�$*E��Mx�C$�=Օ�O�E�.�ygh��
����	��2:��qvx�ۛ
��s����!�u�h?)�Xg�A���I(�XA�e�5<���M�Ȓ�UAw�����)&�������R!��!6X���b<�f�hU��,�'<�1&��,>��<�<�L�`,�d���B�1 j�3Z�V#�W8�<zBB�����I��&4~3N�S`�nlYGtJb���Ρ<�K�R��y��F�~�b���A�����.�L��7)��׊�^�hKЇ����`�N�*-w�ux}�rɦ��$0��g�:?���`��
��f�4������D��}"��i�Tp���ֱ.��_K�,�y���>��\R�K�.�J����3I���}��ng!Z-��<V���I�1�[g���u����H�L�}Cqǌ{�h�"��$�����t��K�I�yr�9b)��BHM����ZW�z��_�0Kx�U��^:�+~�-j�@6�9���h�]�$�6쬍Ԯs�C��$�ۀŴ�7�\�|y�"(
���@�bf/LF4�V�f�:��W���xer������K��LZ�� �?^���8�ؕ��T{!4�_
��f�pPGo�W�j.R/9�}A L���b�4K����)��_d�J�E��F�t,��B�m�z"�!�&�i3N�\������7���.I�L�1>���(�7���ַ�<���°O)�(zL
�g#Xg�n�}���Ǌ0�����g	���S(��I�KDH� ��8���G��洒�O*��Ft?�/P��~˞-��E>shq�҄!��TM���?���Z�aɴMK������I�����l��u1��S+B�E��R|	��m�PG��#-��LT�0z~g���qԍ�w�J< D�f�=����We�ܤ3ծ�x˽t�]?C-w�����\���*��w؞b<�E㜓������v��QBO۶8�:��g�dx@���*>6k]Sζ�e]��
 1i�S�� ��}�j�g/	�v$BR��s�x��)���i;L���d`+����Pa���@��@�H"JU�E]�9�v$+�J֭������GU�O�c���X4}���@c�%��r����Q�����}��ZCG�8^��YE�3�/�����(�D=��˜��۾��jԐ�����{�U�"�����ܜ*Æ�TN!�����c{;d��ƈ��������W���ǐc܂�� �N��gBa��)6�(�US�F��\��t�)#w;�4]��3���v�r��<�IH\;�t�g�d��$o��Z�H ��1j�N���G1+�(��p�og�P5����փ �p���&­N�9z~��`�7�Ȍ�JU�F/��k�(�%{i��	H����,�N�N���LƸ��
����%�.��3�R`��l��-"�V�Z��dK�}Xl�թ��v��ؗ�1B���.~�Hk�k��p�i��_l!�f�
���<Z���!�%s�E!���3���C iQhՄ��Ӻa�%T�hEҀ<�mwg /Tsm��X�](���'튢Y��w�)��TS�Ffq�+��dYme]/�@o�y�k�PS�1;<�����J+[-T��X鑠�=R� H��!>V6����+p�,F�~�L�A~�cĶ00�6K��	��|W.�^���
�Q �~��H�8��д�Θ��������I� k��Ó_�|y����I�R�A���9
#܌�$pg����l/�%��)�%��a�^���e��R��]u�ݍ�"̶���ƭ/��ӆ^N2�.�I��epҳ'*�ϼ�>�����(��"`�$^�����W"�IӸ4�k�#_�=qW꠨;�nN�=� ���f�wr@�ח2YII�o�~mIʍ�u�t����XA_����1��L~�ɬ}ӓ1��½����P������@�.:���l�ƉpX����-����aE�^*��5c�� �77H-?��S)�����}���n�%����n_A��n�i#�v15:nV�<Mx�s���b��3.V�L�00�����"9iq���ƥ�l�8���wG*��v��9~��
�YX͙G�m�]j�t�Ǻ�;yt0��̈́�us/kT�-�_��D�~Mg��4\�F����*�DB�G���#�	z!=q�>��mMغ��7��잠��C���rG�������/�!�`��UM6+fg���wx��E�M���)�Sa:�iJ���4�{���v�������/�[�qHW�0GO�r!���N�����ƺMTDܢ�>�����xQȩݷ�@��Zx����m�����dv�ő	��ė��=<��m&h� j>Yv4!�)�S�~-҉LN+Ť8��B@rb�32@D7�S��%��-ᥪ��j8%'!+/�SʂJJ��-�څ�P���F���'���[2b�m����,	^S�JgJ��2��{�Ps������s�B�.�~8n���~�#)g�bYZ���"/V�.���?��؏~�Dlumu�]�@<�q�r�1�2�e���`x�����̺�w �3|�<�r�@f	\��
�YO�A�@�~fC"�a�ȇ��K㱟�nᕲ7Z�M�t�x?hGC�Lq�V�.��h��)��(�y���:��r��p�yǹ�T;7�l�>*�D�7z���W���H�g�6>�G���f���`9Z��|�{vĉڇ(1��+�˾^ogt�p͢�:���(���h���`�gt� z�K���v9ԫ���S~���,��������P���!�E�Uyl��-s���wV_��Ŷ�5�YS�{�u��mѿ�'��_|�0���̨�`�f���\UO�5��JU 13�L����c| ��im^�l�.%uC�F7�K��Սx`6���u�t���Bv�"�ߢ������nF#~M�s�}�ճ�ă8���H`�-�i�0�а���u�{h���]q�2=M��ŗVK�+���F�R,k�i]�,#J!w������UxG�h��a0���9��rs��D�N��64�ٱ� X�8�И1H7�|��t|�\��i?E�M�T˔ı�{I���� -��&A��4	����k t�.�ɬ7�QO������_�~wu���L���zF(��0���v�}\6Gx$�$Vf(M�"4�FJ���{�P+�(}nb���PǋBTFJ������/�;wU1�Lm�/�M������I�Q����h�7p�3��c;uc_w|% �=���I:X�/������/�j	O���x�C=��m��������2W(P̼g���+�@*��D@ 7�U,�t{����\�W9U�J9�����J�'O��Cj�Ӂ+X�Ϟ�x��� �~8�aԼw;�� �a;wi��mb�D��<<& e�P�y>��7-�`x#���#ȩ�����Iz ��0�h��%O�۫�|ĜA�����DX�X/6�Ҏ�57������ir��Jx PQ8~�w`��&�F�����Jj~�8YJ�Z�F(^`�,Կ�-���~A�/�j`/D�"�Fa'��X�r�b&;�<)��ߑR����Uau� c{�Y<:w��̩?��x"'�Fw2��o��``m�����Zh�G!1�)�ÊR;Xzu\�]�X��n���DUUa���!��u�pw�������"]U�2���%Gst��Pc �d��r"�,���P���gC7���� ��ڐ4	��ʘ�C� �I/�B�IG�����Q@�8!!K!��K�[O1U���)����B�BK��e�ZZ%�n��U;$Z�hJ�/�{YB�밌c9lc�4��@Zz�*a{�ؑi�i�u`�c�(�w�0�E���`m�-����<W8�ݗnҔ��2�i[q��H�J?%��Ca��R�ȧA�h���Y�D� v@QOP���;��TJKU�gO�-2pv�\<�9����
�-��w���^8M�c���>�6��iÏK�f����Q����p�;�o�xF�����c�5:��4�(���Ya�L�B������@O���o9�x�]��쀡��$�F��;^Z6@l���$��n��cJj._�@Ʀlݸ	T`�0�<��������ת?q���U(t��H"�3U��;W�������v��Ħ���\��H�K"^ ԿoF�#\N���k��Q ��GYX�,���쮑�%�^r�����qK�� ��6��Mr����ҋ"!o��sى�q�N�[d�`d\�4�5g"6�w|������xN�_�&:��Jd���������w��yX3�e�7���	}�v����h
tTCr�	��/��޶�n�s��sqK�0
�|���u��7�A�L���1��*��$��p�G������Z�/���s�'�%�!_P]O���lĥFW�����w9u����b�>���7�k����l��r2b�u��T?WE�|��kԡ5�tE���jh,��������_���^�P9�g�MN�4H���9���s�^�H�ăަ�,4]X�n�2�l�aw�UlZ�R��I;�#Q`9طň��=���r�Ew� ���oI-�I��ObY�z���ɞU2e�R��Kt�S?te��l<mX��4�0S��2D^��h����N�$ѩ�6>E�Q���oe���J�����N���p��L+J���tge�B�B�.X�Yl"j�ǌ���:��3ð ���_�L� ��8B�����r$�I��	��V�6��(���G�ɂ����n�]�n�p���h	�Ӝ�6q��m5�ĂE����l�B*�j��E솅�y P�d���U����QKC���}����Ys�B�j*[����؟I�ACz`b�A�=�ae�7��?�~�;c��j�Ú.v
�V)�o��N�X}T<6��'�G0�ݧ�Qup��
a���)�_�Or�XlxVHYEB    fa00    1600�bx�&�Ң� �mk0о7N1��BV:��!f�\�U����j�tZB��huG�s�g���ٵ�Q�GL�2�/h��.�d7s��YI���Ew�F-�,i�����L�OJ�]
���Üs;�fZӖ�4G6|�A�}�0M�*>�2pA}&�K���'C=L��D|�&kcc%]Zx� ����q/�t����#���'m����M��x�'��(��2@E��J���ڭh7l��Û5�)#�wO��/5�U2��{�K
��l�cX@�}�\�,��8�]&1P��t��w��Xj�P����P��H}�)o*�/�J:���_[Y�S��o�%t@R*زv0��C����l�]�t���+؃O%D���!�R^�qCO�W��v�R��D�>���FU����U�������*�C��cu@B�� �(L���7�,ͮ����8�!�C�8M)#�z�� ��r�b`�j��l����"��r0$2����)Y�,�2�b�ck�ą{|gxTC)w����~g��)gj���Lq�Q�G�Jf0v���2�J��dǪ�����N�򶎗��x��=�_��>�W$ɾ�g���,m	�0�����
&�Zf�ç�/�A�lٯ5�9F7e_|{� ��)����Q|`�l�^�2�N�WvʙJ..y���|j���E��"����L�=��?���_�%3�~oi���Cp��t�FGw�c+0#�,C��L�L���\,���=���ױ!]��'����?�"��u��KP[�H��@��D�om;v�����2�%7d	���\~ S'��D:���ˮ��b�)Ҽ0�r�E{��oؑ{�^�r�C?V~h��;ˎ"xl�j{�\�R��"�u��[�i�»z�ao�0p�H�Y4%���pQ�+���2S�����栆���R�A<
����D����坽�/M�[f��?Ѻ�ZϴM����nj���t�-������W�&���&����#��[�j%)��!V�[�[���:J�y;�����Gb�x�e��_����#���Z���zFZ��3�v<��л�З��tcׇ�Z�1rJ�E���.	ܛWn�+�	�����Ǡ5�]�����k�`��֛#���f$'��v�i��QZ��@h'�	�l*�ҠE��%zx8x�12ɶ·1�<�aR9{C����k��j����qDP��J\Y�u�>�J��P#�/���.�$��i�in�cU�ƓZ��"%I��uCn۹�FF����咫{��@�a�f�Ϧ��Y�Z��n�J9@H���a]D7���D�y^��p�\����6�T��<f�Z	�B=��:4��+����j1ݔ�P�q
_&g����y�Xp��-��~��H�P��C����\�ʩg����m�԰S�9��U�a7O !�Mf㑯hH���D�(��\��5V��{�I���Z66�a��Is��miIm�2 ���zF)n�K:P�i���H���O�ыlG_mR�*}$�ˎ|��W{u�����?��!\�EϽ�7��Ӽ1km��+8A�����|��1�qvaAQ�%��B�8�iA龈jԭ�C�$�6�Y���
j�k�!V�c�x
�A�7f��\�ŢO7���NM��@X�@��:��k��^�	��['��\B$n�U�T�Ԝd݁>bt�wN���@�u�(nv��y�{��Lv���G��I�ú@>�<m�,�E΄^Ѝs$e)I���o{7��m���\��%��w�;��늛�h�8R�f�K�5���/�z��CTJ�Fh�Ų�간ܱ������+elA1i�lM���}���w@�s�4Ճ3S���.*Bsc&�h�z����}���A�2R� zӟ�1�8���- �ᬮ��O����FT:n�#�~��X�6�g����Ьc���x�pҮ���گ�a
ͥ���3ͮ	<�;S'D4��W-\0��G�P���;�w7�!IB*�1�N����aj.�CR�\y�o!N����*���t�\LDvz�Քi�M��/���<�ޭ53[�t+^���_.WvZ7���ib��cC�J�"9��Q�SB��,T���$^Vb!^���	��)K��n(������bĊ�m���j�mM��"tG �I�x"�Ѡ��u�K�կ�q)
���#�������-�l��6J�A������\�y�TwG�6�j8ۆK0�˙�A?���x��|�U��E�!9;2�E��v6L�x��]���d�/ƚ/��2=��ڢi���.�AGrZy����9q��m�J��.����0��F?o|i�{7gj��}�S��5U���`�^�	��϶�����T>k�-��<�@�ȵ��Z��E��"FuՍǃ�*!zQ�qT���F�W��3z��8{�3��`�����=��Q�P�c�%�$���?�B�@�;���F�=$c�J+k��c �)�7�_��ܓ���O��W{���?6-V� $�s&*���v��u����r�^��>�
)���"��l1x�*{���».����!�u�j���������3�R�ᥛMz��e Tn�[��dF���@8�nd:��F-?V�e��SΠ���(!��R��Y��W-G��� �����1ty���r��PͷO�PT�`_�j�(�aU/�;�9�`���2�zRd:!�̌�D���g�x	�[P	n��s�"y���k���p���L�w���l.R��r��T���3DO�!g�W�̷gǴy��t���Q��:xNvE�� +���D����$}FF���Y���z�N����Nwq��U�`Z,E?U��蛖ulfDVL���)?
��ܨ7���om�[k�R��	g��^���[�m1y�Y����-"��ݶ�x�8��g��"9X��O*I��  j���_Ώwlw��	C�r�W�C���\x)�z?U�Y�x�E��9K]mCL\�d�f��`Ș����d��,Ձ
&�5+�@��6�m�$lui�Ð��1y��8r�G�z3W���_V���(o���a�9hPK�����dP���0#�	�|<�ͫ��q'�O-;�U��s����Qy:�O5�@��ڨ�*�^��:�����b����Y�#4T>G���ҁ}����fΤ����˫9���[��*d�/V�#2�.��1�#�.m	7� ���Z!��_#���g�R����M�a�J�D�G?K.��	bM�[q<ڐ�s����ORâR��K��n8���	\��H �t�4{ZӉ��յ�Dm�؁爸9X9��Cl[���S��|��7�t��vz�W� �-�!�����!�Ϥ�{�=��T�i�=�d�Nd��tU�)ݥ���.��,���t�H��|��c�+��e�J��� ������h��5P��w�M��1��$	XC���8ߵ�4�tىЦVz���&
u��}#n�.��/�ے������5�_�}�
�2R0)�F�v�B�~[(�K��m#� �o�?yJ�,���_\$m^�6uU2�R���MO�+�iҦ���6`޼^Ao���_2��1/�ʗ�;.�}+0�6���2u����}
Rh��M�.�Fg�s[du��$��C���p��B�o0���-�MY2��6�{w�`W���-
ND}<����%��w>�?A�x{t�c^�^��<�사�x
��ũgZ��aS��M�H'�F(�2�ly��<ސ{Xm��8�LS��\��c�^�k3�Y%�čP�8b��pE��[��aa3Q)�ًh�4&��sZ��GUʹ:E�(k�ޓ1Q�zm�sA��m<U�k�������m�{��S��bQV����NH��w�lyU���Gh���i����יJ�=�}[n!�K�jS�ߒ-�퟈8��2ԑ0�X��y4�RD�H;��I(V�!�g��M�����9D��;�I��j�©����煮3YX��W���$g� 87�_�+�7E�q��p9%���^423:#��
¦�|�k���A�Ed�)���5D���sC��r�4�'���پ�ȩW��	�{A�MU�7�pr.;BҞ�h�3j:��\�T��>h�Ő��@,�f��X�enp��s�Y�j�2����.(T�|u�B�3,�ny"�B�?=#�͡(���-��<�7O��_|��Sl�K�xl}�¹g���ȸ����+6���B���`b�Fi��Ai��]a���X�$b��\A�\����oL�F��g������Y�X�>��]��G<m&`�!枽:������*o�S�y���N���M��9BYηz�g�u�� E���e�&�$��Ϗ�7{UJ�K�1[�B}��v���VF���s��w�k��`sZP��9�#*%	��R��Ad����H��?6��Q\�Ȃ%M�S���8,�.e"@j�bN5R򬩈��� �A6���_L@)2~ChB�t����%���F4�TG4��ܭpPRI�/�_ć��K�m�S����	���(=��*�n=T-� �_m?��1��+c�&���*��ߦԐ��J�۰~'�t2wX��.� �a3��Ǡ����XZ�A����ܙJ�mMr�@LV���ѥo�=SX)L+j[U������n�V=L�����A$�!͗U�ET��N<�ƕ�%��L�F�3�Uqj�����wн��V��F���	�Z�C��ρ�˩義~�[�O�`�Ű��L���ˎu�����F�i]� 4�3	�g����}{?US�����6G�'����GC~�/s�1��u��Q� e���"��JN���6�D��H]�x�s'޻<��~���G�I�V�M�Q��B��K0;�����(��m#M:*��w�J�u�'� 㫂M��C��#0[㮜��^�T��XA����U�����^�O7�|{	�w6��d{n�\�k�oJ���mG*�͕�hN����-�T2��7��H��R6�LX��j�P��~s*���.g�j��.��_2��@MGp��u	�z�ۍG���{���,��D�ctR��6��qB����=>� V��I�-W0����ݑ5Fb�T�e�=�;}~ہ1�0s��|���Z� �;�;VjJ�:��!���M,�O��"һ�O5J���]��Jd�ff:�{8�c�ʾ�Hr1'�O������P(���]?���~�Z��8�*k�i6ߠN�J���u�?��I�=���]�#T^��3��QQun�DZD��8*b�
[��9ev�6x��[��NR�W���mS��Fa�*l����7f}�i����1�b��c�	�0[��P��j��0ٶ&���U6��B��ǣ'ԭ��V]ˀkB �J����㬼���ZxO��qV�M%79�ce���vk�X��H����_N��w���àr褓�Y`���d��;�l��im,l$���魜
Fj;���Il4���T�N�)dv9��N�ߠ,J2���Շ�:�H�E�,�l�P�=���m�=��0��̶��˅�XlxVHYEB    fa00    16303(Ԣ2>V��BbH�b�A�
�-��]S�Yg.�r/����E��<��U(�/��pVI��R@}�_��=���aW[�'na�\Pe��Ix��aN{��wW�_��S�!��s�:B2�6Ա3
2��}����	�����Ⱥ�La8���]�a�om�/r���Kn�(���c�����[?�����#ݔ�6��@��!׌������� tO��iP�
��|���noק����C�uB�:;.��wW�0ĻY�6w����f�P����6�Rpj�Z�i�S�r��S׸ �n�;�i�rU<�:4�ۭ��_�x��N#N�9i<�������9�4! �er9ՔsZ�����5��f2���㉩K�0䘿���B��+>%=�	�<CK*�-f.z�:���D�X=DZ�L�XY�?�;�Փ|��J�cf@kI�Z�$A�9b��q=�rPp�3��&#ȂM�$��\�yEqI�(LP��E���p+k#��"��gu�df(PD���Q--�ь1�*7�k��k=2�0�'��P���]C�_�p[bO�2�C5�c�-����O6\!�X7�!�\_lg�C������-���x�_QUdM�$�
o�x�#�a\�%[8}ߔ��L�-Z^-ݔ���~�.�����u��(���Sr��A�S��_�<��l?����-��.�g��Q�W,~v�{�pXhB�����gζ�~<>J��k|*�s|T�F�,`(D޵2���������yc��cS6r�.�u�w���5nM���E�,vV�ھ�U����r�UYG����]��f��I�y��Yv�7� ����34�V ����F��]; E�h3��'��,>�b|�*S������\��ĨE��܁3
����A��x�t�(aƧ+43"�v�'�B��qlI��[I���,AG*�
[�M�����1��-�Iٕ�]�rguU��zr\����S�YGۤ�k�K��&Cf:�ܗ�˂F�������u��n�Y��H�'Ģdҳ�ߡ�u���i��t���7��*i���q���f���=H4�e�L)�_� �Ͳ��:��zF����굽2��V�F��g��17x	�}ER�W�k���M�F��B��6�#�WW���`��|����Mh����jW��R8��e����a�����+�	�"���7ɿ)ߝT?�A�X��#rg����zq�*$� ^*�]1�Q��Gb�Ijv2�ʙ���6#1JDq�B;Эܦ�P�B��o�١DS�:Q��s�W����Z}����z��1d�:�ۢ}/��������S H���[��QU"3�'n����b�IK�xD�����E�%�d�{�8`�Z�G��+Z�N�cq!&F3`i�th��˒��lO� ���?��]c�t9����֐�=|wG7�Í��T���=K�>�?q�9}@�*?U�!�yř2��AW+����p�ο9��7��#,!>���]����(��tp2�"�̷�M�(I��}w��[��f�)��<!R R�K3x)�~�
+B������)E՘�KA�0I}F��\i�!AʺaL_s��[�8�j0�������T��l�����"aZͬ
�W0q�� �kGB_����|�!V�4Ơ�ݹ�Y����MLΫS@,f��[���'g+�(КE���Ȓ�P�پ�>�T\۫� ,��X�	Y�Ҳי�ߥڎ:]�!�q����;���� ��X�'y��܍`EL�{����)Z� w��@����i�&`����mg>��ad��-���ʻ`��a��ې��d[����}�7����2��v;O��6�g�F���=�� C�2�Q���쿔q���=�^� �KQ������Ç�u5E��#���r�;˷c��ݱX;�>��|�lT�ƛ�������-6"�z�cp�ƙ+���8��3<0��w��UjF��]7�H~3q1^��W�Ή^ř�шP�b�O��1w�O�I'����w��Hz(A�[а9ݦ��)VaGޮ�s \��n�%`ٻm;Sd�-�R�-V�㼩�M�8�����+�ݘS�����4O��2p[�!G�j8X<r^�Z�L)ᘚ�}G��%��@:N��Qnw@~h6���D5�kci�3�A5�H��˦b��S�0��s�kR<���z��Y6j- �VYε"�m��Ў�����))2�)z$��ڈn�^��k<�?O�޴~�I�M���"�|�6M�a���`����$���^Ԉ8*��T��ˮ52�=I���i�)'	u�^�d�4�Ó����ʢ�˙]|y������l�;�ot)�M��8��|�_־�<�_F~�~�Pݳ�L(]q)���`3�M�iMC;��\?�Sܫ�Ӡt��Hg��n��mrSR���y?^E"c�5V�S�+�B�9�;���M�N;�j��P.�`?~6{DƵ�#v#��YP왲]�.�R7�X2�'�e��w�[�R�,���VЈ�����U_D���U
�E�M� ��\�1;wK�ԝ�2/�g1��CnM6\f��+��	7�q1���u�ԍ�"~8�����?Yj�� �M��J7c�K}�Y��>AHl��ӎ��E8fi��
 �Ҿ��� ��%/��̔{����@��]�l(�q��&��pm�4�}U�U�����ݟ_��)i�c��}����p��o$�W�_&��B
�O7K)D'��|���Q��:>*�h~<{�hS
d�E�d�^{hb�A�+#��ÄY�;S��o�মM�M�+;`�z� ��!��"K��������b2��oN�B�,B6���6��m�B�o4�.��A r-�I����u���lֶ��942��3�JFCr"���&P�9 Á��y�>]�k	J�-̓H|W������ ��6�i�	��!?c:c誖8a�����)���::�-�Y=������˛�ߊ�����^W���H@P@��I��J8QDջ�	�P��g�?��]�wf0��E.�E�.�aCd!�*ρ��B܍����.`F3V��H�V��y����ɽ���D�����4a����9p�d�G`�p߬��U@V�h�`��Q��{�����56G���-Vg�[�U�`;�����R���Ek½sY� �[���:�#|��އL��G�Z��$� w	TO)P7�����q9$�g䉸7��_$���2	V��f<G*���(d�urH�J2S@��b��|@聄�]�a`��<p\����"/�����:+��6H)��J�3΄S���5pP��"��52e��p�U�Yc�>,���ڙ,G�l�q�7�l#ё��K�lk�eaaK,���L�*R�����E���:��ı9g�}�$}&k��t�,�(3�2��a��L�R�p긼���>r���N&H>ra�^����g�U�����P�_���|:X�p�V���z���%�ǀ�ӽr�U��.�N7�%o�?��u�Ӭ�;��{Gs�
�K��5x6�"C��Z!��v�x����dd��M�!��r�ˈ�<PT�U��N�߰@�'Ll�R��ڠ%��c��j%E��_�S��%^���Vs/ýq$��X����dn�X,up=��!��}������V�8�jN�v 8CIg����>�˳�PT����J��P{�r7��&�"���=��0��~+��|���un0W�:�끛�w+0M���(2Η?c}������b� >�~��"���xx��'z~�Mj��+uK�`���M�q��*�]����#󅐁s���R�aZ%1w�����2):hT�̋K�"U?�fF�y@@
���>4��R�U���"���<_J%Κ)ݶ��Q�J���� Q�B��@�T�,��g�pb*r��m�Pٛ��#i~ư�y���J��rP4�|-$�%�@�Y��\��Vt�M��~���s�����"�r�6Ś-w���7�gբZ}M/0$B������ȸ.bWߴ3r�b:'�ay��z�}�͊�%��M�'�A,P;io|���q荦�:�H!��S̩;���j;~_�1Ec(��;ջ5�]X���y���I4R�N�m����;K�?�k�y?ټ�P�����H�[L�y'}jL�w��w/�j`���j�O�\�K21#���Cbj��\i�"eI��)�z�w�O�-r�ed2_�Bh�O�O����\e�uw8�$a��A�m���*�n�)?M�Ub�$�XKjej��}�
���;O���S�&����sM< �[���8a�j�`%wl]��ǲ���(k6����0�vP�a�`	Y@?p8�ۥ4a_3Z�d�	q��6
�}<��6�AMQ:��*�u��g̔��\��	� �5�%U���H�j@@9K�<��bë��$+Nܲk�F�i;af�fD���>���Rq����&�23M�;���#��M��t�ɬ����}{,Uz�i��͢�H��.��i\�ؒ-~��~1���NO`Pa���mN]j��U!��UyGd�����v}<��P&��܎u�r�*&.���1ۗ���p�I0e�ʑ����<�=}���+~�׶y������tXɓu_�I��1c��o�X:y��V:�)��� ^���� c>�Er�t��6Fe�1lA�N���<���Nւ�}nP���~�CZR�����?�+�$7{x���a*������<=�>��cv>
����D`rr~6����	X4�;E�,�_M3oQ~���Loں[��r%�oIr�3���6'�;���%٥stcнR�kj�<$W0'o@�ʪ������M�T���q�v�6"ہUC��2��O�&�P��.|��4;�d���P�Q6�a�"���`x8��4�$�q��� ���n[垌Z���XSi��Jt �LN��23�''�4���ť�Nn�A�������}Z�Ņ�y��倨��3�]��aJ��aY��A���Q�mA�d�CYge�cU��Kg��U��M˔r�S,������#��+�s���S]ĸ��Ȯ�����ܰ��M���"��F��;~f��&�\(�J~�i�N�#祸,=|)�`2`,o�;�
�04�j�8�i��<1�\O��#?���G�:�^)r�������]�J�����}\��7�>�l�B13G&uz�������jt�bkl���M˻ss%߿�`�����b��\�c�� ��i����'�|&L!w�u~�hC(��l!rR�-�u��tr��y����I�W� �% AؓW��i1��E8�߽a�і�{�o�*��(��0eg�~�20{�KXJw�NS*;�P|5����R�Dh.u��v�$�7�[E��*u_�agKyB���=�l覌���r�1�H����g�:�#�0D�1��k�o�P]�&_��r/�U��w>�<AX�N��v_�/a�76ho��2\jM�e������Rc	�!e�?v�|���U1�U�g�s��cXAؖЉwb\�[
L�M:?J��i`<�֧Y�v�xX���l��|%u�Z�n�ۦ�Q���.|�e� ��XlxVHYEB    fa00    1620�R��U�ړ_E��J�4�n1b����BHN��kC\�	GsKh�?\SL���.��~쇏k���
�ޓ�~��l�����?�I�S��57��5��Ǌ|oUy�uZh��'���R��0�8d
*�x�B�RdGh�>t�I��yE�Y�2Z-^k�@w�<� �M�D��H@{#�`����*�i떅h�v��N�e8Z�`�54�U��
G���(�8	In4V�X���Gh���}G�+M�����UeM���TD0�t��*��'��'b�O���$����$e,h��Gw�2�����4�	�͕3%̴���ƺگ�QDD�;e��`3Uh�lQ��R�wf��I
n[Nh��B}��h��ݬ����HM����z"��Gi����I޹"��pEYo��44g|������l�W5l'����+&����z��x ū��������ec��m2}���47:�Gu�o����@����hlO58H*���{!��wI�KBnWԚ�λ�'��>,�o ��c�ԃ�_���ͳ��8;���O���<%׬7m�t�Ɗ��;J3���o}%�s٠�xX�ݦ�z�AM��(��R���l�b	
r���^ Q� �4l��Ռ�������F8�{�>u�4�4�77�����]�9Й8.�۝MU�e�&H��N�q�Q]��N��/Rb�6���ee���kG'Z�h|�`T���Ȱ�=�O����:{��I��O�����,|T&�C:CV���)�Eɿ	�(׀(I�ζ�'�$/3p8|�|kl���h�]�8:���2��fL���7e*%+jfɠqs�ț����ꥂ�ڣ3�0?����kl���4,��@�}�;p�A�	�TX'r���tf�~ȶ;L	����q�yIt��ac�,��
�ė�cȻ4�s�1��џ�uBa�m�0�G]W�����aX�5�&}?3���ʫ-Z��9֜�V�Z�B�f�q�}Ew A�抱y��=������uE�ф�IW�����!O�G�۵�҃l��-E9�>����k��W�%&�*H�*G��ym	#���`��d�)��D��{�;~�QM���
��`M0����Ψ�J��z�P��<e�OCw.v����]�y����,�m��bƛ��UZ속ۤu�� KB����l�_u]�¸Si8��Oʋn��ZXV�k9�o&�]��N�́Og��ϓf��@�hu1�HPH�jN"���2�Z!��������G�T��ª��8� �a�����a��!h��v>}�o�ƣ��ڲQ���
)�T[����yۄ����/'�S�� ���gcR,�lq�M-��o�--����~�y�ŗp1L����sF�X����_�\txbY���%`����+6���++�:Io��3F ����%�+�sԗw©h"��,`y+]�X��ѣ�ݛ���"���R���O�Y#�fNfw�7VR��U=�)��ah��mӗO$�	p�eiK��b��^ V�j��1�����Vg;ܾ�ċ~�`�̦肋���/�-�W��/T����R������N]��-�Ť�u���޽��j��`�so����j��g�:՘�Ȯ�^ݖ��m��x 2��.��ۻ�`j��	&Y�v�P(c��fq��@�c�R�rͫ�+�k�G��j}&F{���>�ofr�=}g�m�l�q祖Y��c�3���A��a��s�*�u�<�������JQ�t�T��Sq��?aMn���f�H��6��Lg�3��̜?6[�/.��}�*���R<NN��(���E��8~Ŷ"��/w�H�{^?!�3;�Q#��m8Q��&�p@ʘ���� a3�W�I	����\Z��W�uk�q y��1&'�*�ջ���'g�Y�Ģu!{l�p�%��q�u�]c�`��q.�1֝��pDm�cB���Z"��c~4����[;j 4~��I8u3��|'[b��8Ҁ�;[��<_���6[:��0<�'M6E��'��xa��=�
3ӡ�{q�R�3n�]����o�xR����Thh���}v]m�� ����]����J����H��o�S�����STG���s����� !?{��}�(�4�yЇښ�ݻ�!���e�0���&�%^���&J�Ú����?jc�4N�G�����
���R�X�t�H�)�!YWJPu��NRw<���]ַ�}VR^���#U��>��J�ˁ��8����l��Q����B�Zy��%mM��O���9}C��_�j�l=��> �"A�LPsL�U���4�!�Y#���=n	^�����
[�f�2/g8�Қ���zf�7O���xM[Zω΅.Y���m�"!�B�����D��n'E�mNa�v���}ʭ�d�cLFc2��0�ϐ��L#�#�Ot�(�a��f!J��osw6�'�1����օ��A�R�9�V�g�btѭ�����2�s=s>����z�# ��ǖ�a_?ݡ��)Tً�z���\>'��	��|�/�v�F�w�l�h�+��}�ԋ��Fl�q��P��-�i5i:q�f ���n���q�n6�]o�����2v;�O<�����zz�5�X��wv��'])����}�ؑ6K>��d�t;f'4�]���_#%!��y�ǝy}@i:}$i�����A��qE��N�)�=O3>Jx>r�I���	ﯳ����~~���M��ߏ�H���mF��C��@a��0�}�t�Q�N�"�(x�1���WR�Y�I~�ta�	2������Х1~�(�W�&��=ǖB}�q��i�3�U�N�;\�=*W_�IYH�>y��Ƣ�l�a�X�a>b�����S8�f����J��+�4�*Ì/����l���B�K�!�V;�rک�:�*���$�a~���/5I��@�AF���&�T¨��|暠��}�ip��
�U����"�<D��E�W���]���؃��$��H�Y���i�n�ۄAT�i�4U��BO��sf�_���5 ���~ی"�V���>�ɻ ��KR^]�F�(���c����@-Y�J��#/�J>^n�f#�k/���"�3S��믂��,����ZY�[o��C0�9<�}w~�d�	�!�D%.�{I�j�zH��#���^����y~T�q���4d�8�+A�s����� �R$J�~�}~u��I��}��gK���^��e�KL*}��HU$����#!8V�mu�ob흉�u�-�w:�:a�VwY�r�+��R��0�ů�*}��	U/I8҉R?8�>IǾ�T�\�: wvo�BJ�V�6�IBz3*_�C!X���Q<�1�/+ܑ~�V|����8x<�~=qT����΅Ԑn�G��t�Q?S��e}jɾI�%���&=	�x3�r�.�>�� c���'�f؊�	!�Rw�>ְ�:�%>Hu�U�φ��ĐT���a�>�ʃ���Y��o��?�Cq�?� ��}�,�m.o85���K^(���� �K-S��jƤ
F,b	'�u@��M�qu�	ěk!��D4�ɽ�0�myG���d��Y��R^b����X�(��^�ߩ'��3��ߎ��{���3��h9��vD[���BcG*����6f�#e�&�m���c�7�=U�jQ{�?H�D�P�U��y���(��ޑ�'�8��Ĕw7���ج�kt�Ƞ�B������_\�~�>%�5�Z����R�����=��&�ʌ�<�pEr0�L웑��-Ћ��ݘU~���ֽ�k���Ԩ!!�&�Ľa~N�S��Rfcr���pA���#��~�?ٸrk������v��5��`��d�͞5����9�e3�>(%��,�GWF�=܉�:�6�#�~�����?�Zz��}�I�<M<�#=��Grp�j5�<)o�iD�l�8�N尔)°�zd�#P�*h(y������mω��ToK�*���J��n=�j�d��Y��duCU���h�*�6E��a���m@��@o�$Uj,;JU���[�>U-"1gܘk �����1��N)`����Q	%�%V>�G�i� ����9U���PJM�d*���N|n��Mh=���u�ADVB��)z=b���+5m͟�n	��'/YF��)|�x�N6�P*u�1�.��$�ZR#P#�k��Ʀ����e֟����L��t�S�w)o\�p���N�]&��3��/rL�ytC�o�+a>�P�)���N�U���dԖ��问���t��3^�)�y�;��YK���Gp���5#�<���"ӖR�f_����㵏k���$��k��Y�;�Ӹ��Ȧ~4^B�Eɝ������)M��K���m��<U|�8zSq��LM'���%����iwj5�ϵ$�J۩�N��'��za>�G�H��i]�W��d�Ek����7��R7�7n��x�J���9ʇY����l��5�rN��0R���t�g� �w��by�vG���L�9ũ����8gQ��N�ĵ?�y�l�9��WcR�}�t�rE��X�2�.�т��	ҽ� �:̤'���7����KW4"��E�?���|�Ze�ɂw���N��9i��4�]��\�����ǐM
�o��@Ry4�W�b��x�IV߉�X4Rn��̓IM�s�O��	"KlX���ߠ��ǈ��HJ^DE�i k���em.an���R�i�hezd��"�3�[w8 ����3����x�V������>��9.�_BФ`�@%?�;/P��@q���{E�(Y�!w�)�ueK�(�6���Ƨ���ay'�=�)/6��l�4��2�^��g�˚0�;�pܖ!%N7>ʝ��J�����N�?�����x��M~�	�	ʒ��~}n��z��1Q���Q顎��6Z'��Ϲ��-�9�Go]�����ե�Pd�{����.1���5�����0�rр����̢�X��iU=�=K�i�fo�	>J;oT�W�ص�e�{����w�m]���Š���}�3
�=�[U:�yX����fJ�}Ö9�y�Лh]sO;���<�r�]I�=
j�W�m�����(�$�Nl�Ώ30?��<C 1F3n��.onbi1J�·#"��m�|�诖�{h)�����!���G�jp��;o'7	��X%D{wJKͼ��$�ϻ"�����5O����0�3��2C�l�Z�ڈ>�2�b?�!EK������@�ceN���ͽ+�=u������x������[��\�į���eZ���f�Z%����w�i�S0oN@�<��m��<�݀F�`���z>��0�BYu����*��n2�(+7U��U,��G�7-g��}:9��Cy�"Ϻ+6EE�  �7
 �`�e���_X@�C�fO��8�ճ�ft��C����3I��^�R�p 9�RWی[(�px���8}�Ǘ�����m� I!T�QBt�G��nw�Z�V��}P)��<*��W��|)��1�"���t�[���o��6$��>��S��p@�<���Џ���|���v�ٹ=��J)��p l�+���G͘v�I���� 	W1jzC�'ډ�Zra|A��H���XlxVHYEB    fa00    1630ﱾ�̯Q���0�)�A�|��R�@���De�s�O�	L�٤�O�1�ť0�u��?�nMNd�Ɗu�֞\����R
�hy�E���&�+heә��@,�ZJ���(�fWPokF'��y��1&�l�d���%f�����&�(׻���Z<0�*�*)���j<S�a�h<���G��R#����֍�s�\����Ťd7�l"LuU6�aIo��c;��gL����xd�i+�jd�����aĭ&��k�vER ����B�6}���'��Y3)��#0O�n�?�|�e(��H��Z1TV���g�!��Q�ٹww�{)C����K�\Y�~�xA%ց�^r��i�~k�,qC��U7��`��UU����{����u�y@�KzQ��B^kpF�)�g�N�=����~�&���:�)��+
�Ц�Hmw�ҲZ���{9G0~jؗ���}WU�UL(1ӵ�;4� ��B�Z+̕��xG�ߩY�<>G��"z�SL�q �is-��V��"ſ�#�VR��{�'���e.�CO�0���8���C��<U��?��7�����l!�a�n�dp��ݚ��W7���Q0�	,��k06+���a�_(�	�eбJ�@L�����D�h����{��i��u�����ˤ1d��Y`0���P%�D$ �냬 ���J����@�gB�"�R{K�v���g��%���h�fٳ�O��]��eƿ��<GJ���A�(!C�VM+9�?/��!�2}�'.�U�F��ıۨ5�G#XY`���[ѐ.�U):m�Ȩp��kR�~7��~;���t��)d:A[d2�ґ��	Uf@}�F.��r�������t���r��۸�t����go�h�M~0�(���>��J��g{q�V�0W�OpE�)�7���[�9���Y��g�舄6�)�����D� \9��Vgw]�;(�Ro�c�G�H���R �����qW�y%����
ze����v<���N;�Ɲa���1�}��@��(�=�<χ����0Za3��xyx��k�zXF�>�^M�G�?r!�ԝY{���~�N�Ϗ�v� ��������*�g���}Iz����?��;*)0��_鮲�q���q�@���uv�� ��D���=0����q�M0OB���q�a��R�N�o���,=er�����a[�qo�N�~�M�u���~v�y��-h�;�{�fțɂbPk�Z|�d[�S��&0���<b���]>$w���	����_�.F=���yGs�	Eq~� �`WЁ��RNE(0l�cK����:�����X�M>K��q(p��y��L�WF�j QW��f�G5�.(.�Ϳ���6�#^�]y�y�5˦�+<X�ۖ~�~�;=N@��������M�?��W��P�#*j\8qv!AlN{RU�Bv&E|&̀�	���!�wO�)���n�
B&���~�d�9��f�0n���yX��\P�%��im�9,����$z��GO��Vˢc�W��r�|Y(bµ�#�I
�B���&���;X������{_K{�y=re�r�D/H#K�5��Υ�Pߠ ���V�S���"`|���h'� �	jd/Ӈ�<��%a��"Nb%�����h�i����f�
���dr"�f�AopIn;�.{7��\��ڑGZe`�0�����ޝ~�H!?�cYQ��xm���dXH�K�^�]Z󊔢	�/�{�顣�4�.fi�;���4�p�%O6`�����������%�l�|��7N�`��.���ߍ�g(cܵ����)�!�@ŋZ7IC{3D�@�Go�Sr�+��j�� ��@�$)(%���/<�ʧv�*�N*���R�Yb�������X���
���p�kJt�D����T��� ��a3O)l�G��y�M�CÍ����.kX�J*<��,h�𜃅���w6�<�âNQ���w��u��X=q:����=�+o'j�eB��V>4/1�Eh�I0+��������zT�?Q��Z�4r��Yp S���Ȧ�e���+Y?��Z�6E
�\������.�������?/<%��Y��-��e�u���_�>.�q�c�E~ci��Ő�r���m���K�5�'��So�@�z�g1��j�T��Z?H�D0K�O��Z��>Ѿʉ.�Ҥ�I"�Q����1�#�z��|�C)c���9^4J��	hB�}���dƟy(����Gsl��oY��"
QA��[�(-�@�>uR�ؘU��7$����>j��7�����̘�����z^ ��E4*d��U��td�����5W�L_g�P�;B������_n7n�O�?�CB�˂ki;:���<�7%Ds��=:h8�A�t5��s�?�ң�����W��0G�� ;-&� ���~�4�q>��U)��X����1�I�"�+��F콳y	�n�m�F&�j~�ˉ�ze;d �U���xo&W����;3
����Yw>��]=N��&��R!���M�?�zIϮ�d�T��9��]I8���ҽ��iw�]\+HǠ(*!׏�}&�h5}��~T�S�Kz����O��T���������Ni�l�����&��3#�{���F���x�7�}���B8���� y�[����.�ڠ�<�X��|����52�f�ɴ�COS�������R$���xg!�k��G����,ʷ?��{G�BY��,�cm�����1V�7����#���\�Ga���!�r����7P�L��h��<�6���H�n��bއU���,g�����U����E�S:P�0\,��Dl��Ʊɻ���Т�F���g�@Mu�����Y�xXk�������N��kI�.)�Ж�MnK�]��X$1�D����ٺ�/�J�3&���_^�w���9�9��h�0��w//��};Q����(�;�<:yB�7�*G.�vCcU���KJ��9E��i�l�c�4r�&������5�c������d��ә�NU�(�-�n��Y�xXǡ�j�:y���\�3�����s^��]��L)T�~{'�n�~��וJQ���dZ	��w��]wX�߯=]���6w݉$����xRLw,z�nt����s��ON}垠�,��E�n��9��~k+�F����/��#sϚ�;U+h�w�v�!kBB����z�M�c$�z�����FE�7#*���}�o��E�����.PM��m'�2�D��B��3�_�5�m�Q�<7
D^�Ot���e���Ћ�Ϥ��4{���@͓z�}9�`�ȟdݴZc��,�/2����u;�s�č�"��Kѐ�f.���7fK�)ξ�.����{i�wZ�E�O�Ke�����.��&����epu�\g}�a <w=��<�{~�p�?�݆�0K������r*�ֹ�oD�ˢ� :3$�.��N�a��xl-?��X�x�	��K֜���*p�?�(���d������׹_��Tv�
QZw}����o#2��
�MB�JV�ZЃ��� 8%uU����x�p6�����X���K �4/�����p�VB@c���0D�WbTl�D����A;sB�����~�pRv���R.�P)�MnC�����3�d��I��)������p9��N�u0����j��^�&!rzh0D��U�Uy�ѓ�� p���W����\�'��J�qe1�
��;�E6�~�W���� �{s���� �ˇM�}cǄf�SU�����I
�
��u�㑧K*�؞FO���R�mg�\,ί��d�c'���lu��cS�Mg�[��8�=emh�C=ڎwo�<x=1�\j]3�x�B������&ZF3iY݊���}��r����	=���8�q�]���C����{Q��۲�+qEGl�D�_ڝɋ��ɕg��8��uɂ�����E��)�Y�6�Ϊ���o�ܑ����sx
����W�N=��XhL��WB�杁z�+<ˋA�x��V��q�'�7�Ǆ��wLrp#��:�J��f~f�CȌ�M��yjd|�]���!fX =�;~-BlD"�ǜl�\��w��ɺ�w�����D}��M�g�.{wb2��N6�
���W��j�7˱G'L�`q庁b*���JQQ�ܶI�Js8�V�7l�*>�z���[����u�/.�!�)",��3 �J����uq���t�e�S{�x�EҺ$��rk���U=���.�3���u�̨�3F�x��2�ڶP�EgLBQm��Y�J3'b{�w���o�y[��4��괞ą�#��� ���f�t� �3�q5`{�ķ�$�uv�n7�Av)|��Yb�u��?��W�KA��cQ�X5���Z=��+և:�ɐ���Ua	0�aP�E���������?E�Z�~p���'v�b�Ga���$%�����O%̽��Y�D'�(cL�@�a�A�q[qa�u�>�C;X�N��h��X`z���I�8o�]bwr�� ��"v)�������"��\�w�57ݢ��0>�Wa�acOЁ[�&�u/�<d��jp��#���L��Y�S�t�aw���T�C�ϷJ����d� �{���Ց�Q-�����d�XROj����4�� ��U�ZX�4�ڨ	��L�	o`���%�1D#����%/�>��^�,vώ=�j�k��_TZ��Yę�s�}�)Dr��,fbg(9�/��*��sa��+ē���IH���B��s���$NҠ!B�8��6@߰R��1�s���j�@ԑѿ ����hSO��YS�$6�/���"��X��vCTx}JG��q/��'�q�GT%�S���;׏� �w]��z��>��3�#�3��"W���}7�t:�UH��=���]����zw�s�ː#XD�P��#�ϒ˔\��ި�57��%���r��]$�y��g;�$���[s���ծ+R��e���N���1ړ���r��]�4Y�ȶ�C�^�纚��"	D;0%�#�UM.�4[#ݴP��@[X/�7��;\Z>��i1h����3oKz��JF�	M�b]��~ް��+	TNn}�������Ks��8�
I�0�+�[ҫ?Y󚲍WV�`���v���.2LH�<�:�F�]и�MC�׭D�hI�I��1�"#��V�V�!r������6˹������fs�O�{�@�C�!�=�)a�q�Es��jKe�OC�GN8�b��}\���'A��6��IZE��Rű~��%��7pb��5��g9X�@���7�f4�vi���7A���f��r�*��8,��;E���p��q__��^�G����KPcFA��e��TJ���Wi�l�ߴ(����k��s�<��>���kS�4������9L�v�ug�g�:+�9�H*E���k٩t8�C�p��������%�ҷLb"�S�1���Ԁێ��p���ZAV�O�8��ǳ���t�����7���7O���	�ˈ��K{���>�c�]|�oE��i(,HJ��&��������p}��`�h��*�w��%%��q�.�i�t��$5.��j	�D�Q8�\}a�W�ua�$��G�������t�d�����.x�A4{ڲ ��DT�ׄM ��:q��4�XlxVHYEB    5a90     8505&L�.f]�k 28~!�us���c�o���+�Ŭ��ރ�����%��I�ˠ�J秪�n~�dy�V^d��a����!�|�P��0u�B�i�94�t灨���[��w�`��,�^�҄Vܙ48�f�|Q�U�1tJ��+�RQ�>��9�iH߃L�e��zjq%z���Ԅ�;J.�,�Rg��ߵ��������S�2*KN<��-˱\:n��A��-�B�2^�O��-q�n�r������y_���v�^�s����^�����Xd�3,����I�g?j��o�y��|m ���R����B���ܡ�p6��׾L�=t��'�����8G��'���-�^��wɵa	H(�@0��6z�N���v� sc�[�^���h�������%�So�aE����>��=��2eeL�Z#1�x+�����|���:#��V$����2_�l����©J^��䜐��B�˦�㧳	xҚ���^�I#�D�u=�Zw����`қ�k���F͖,v3߼kwҜ{/B�b�H�1���12�-������*�n�2�a�yޣ��E.^I*h-�2��}1�]9Vf���i�!v�b�_�NgUmN��j{-nϤ����WO=��H�EF��2���F�<s�՟xՃl���C�Z���3�x��P1m���]�n�ۓE8�ɟ�=�R b2���EG<�(6e�_��\\3�&$w�����`K�hy]~���~X0<D���L̦� B�	�I�����k�&��Te�:�AoD@|٤����]����Ә�D^ 2��.:9��&�-�{�`�mEM����$��b7�?����t����P6
AQK��)��oͪҘc�I>��V�� j� )S����к��F/{>\w�oD{ڰ�u>�LF����:����r��9" 	��}ʟ9w�U�f�$\�GmK��������͟Xi`�A�Z������HR_��ǀh̒'E�4���z{��©(Gu�	 �,���_	5���V������1�+�A�ay����Q���� ":�<1�n�l$��9�ۏWɽ�u��;=h�'O@漓���ͥrg�=kF�� �l��~�\J�8�[!
��4�9�j/��c��ݛ�*F������E	��1�<��yԦm�u͎���
�cl��O�x�T�(ۑ~U�{�[��4����D}Y��!]��^��b�97D����*߈����}������;F+����y�{�ʻF|�+�xt��G-�eq5�^d�7�����^���}��<�2�x�o���1�P�s�*4�� qQ!GT46P�9�d4^�c
ݧ�gM����x*pq��ﱮ��2ɲ�zB&��P_MA<��Tf��s)kd\����X�К�B?���{s��,��y��L<�_)u�L=����EDWr
�'OO�t��nJ��"��'خ�b�AAt�*F!Ϝy�R|�t�=��z���O}���gn�A)��	�	Dlz}}����zI�̅���^���&q����Hz~�nu���r�F"S�J��|��ز¤��d#�]��
O0���ԇ�J��g4�r����!�9��D)�� �U3	��>�|���]"��'��Z���1��[���,�u�J��1ǟ�$D���y��ʓ�7��&�oc�,L�|���3w�v��S�q	�s��H���PYq�&��@g?'����#2�� ���� ޹��`cdlk,�����%K���2}�m[q��:���Rk	���������X,��k!,!�/�P�4��c���2,���;��d��i�!UM�5D>����J�L�O7�� �Մ���{��x�Fw1�?c\��Kie�7oshS*~~�GG�K ��B��]�'飆T駡I�����h���+�T�����M=��.�A��*��Og�XrJ爡�L�Sꉬ�|=IŠԠ�*7��g�8�������}�['�q#_^g�183	6��V
[�P	�4�p�e�ݫ�X`J����aB9i��
	*)���7�9�_�/�s�x�V����%�(.�蓠�ȇ��GB�v��o.	��Zz@�&�f��/� ����