XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�D@�!����A���,&_�>�c�M�ͤZ]�gq#��X؁�Ԗ	�t�sO�V�����mo�����9x��3��L���q�a��L�-�+��K7-�tX?':��D�/Ge�c�n��$x^��~�]��ц��%��s�_�U���n�_$�z:�':9(����( )/��� *�clLC*t���|Wҟ'�����}�.8~�:��Q΢Q˵b��S��
l2��Փ��,�XYZM�k�5Tg�^�H�U~�8;���=�eepJ���u��G�:��es�u�Q+��d[��WA����}Շs]�y�	�����L��wr��2�h5�Jةk>�a��8�0�����olbyn+X�ɀ��q��/��9���SA�!�`-�cM��2�L��?��Hy�zD�S�)���Z��&�X��o�;tO�[R]^C��a��HJ��7Y��{�Yt�PzJ���[!}�����WAk�����e�:} �SA������Z��?��C%�@]�T�E�.�����~�@I�5:= cI��=�Q�_'6H,���.1u1������K����
)\��=�Lf�O�"D��`��:��jڴf�i�y\Z�m���M�M�$&�ZH2^ٯ-DaD�!��AQb"Νd�qSX�_-H�	O���/\@ANvAox��mz4V��aR�l�6edh��&�Uto�V�UO��2x&�5H@l�ㄼ�K���w�¨2Xy�2�XlxVHYEB    6d0a     be0ev�U-5����_@e�H? %��v��"�҉c�J��Q�܉6q5�2��t�H�����(9���y�m$�mgkv��緯�_^ S��)��h!�<���a��T����.Ok&�XE�E�$���jV�f��9�.�nA�;*1*|�c��AX��\���^��T�&��U��=��0��sT`)����K�����V� �s�GE�VJ������Pyb���u�)��nH�kOǗ���'P�R����b@B}��Zc�}���ϓ�7��U���f��K��1�������مt��L�K�Im� '1��|�x���O��c��b����B����\��{��i7���խ�Y��^N,vg,P�)���e�W=-m+�<�^w��59�Y�"��A���qr �թU���O� m�ؤyŘ�6���g��?o��KGj�f�G	�br��D��/���|c�Ԥ��V8t_�%����	����qg�f��\�"�7����|��n��VI���"N�����D�H�����~�*�S�Dȵ��m�W�ƴ9���� ��L�5Z�SX'���#@�2L���tmt��F�!�̙�m����f�^�m}�� �<����8sDn؟a[bOF��F���د');?���[�t�E;��
��E��'#4T8V� 1���q]�/�
'�7AY�PP�T@'��P���0�؏��؁�Jc~���{N�G=�ܱ�\�JF�PI����Le�D��o�x��6�S�.0G*0�]R��1�u�㯱M��]���潄�VQD6��j�emMHt�����hϳsw��#�7�@������%����H����]@���AF��\��s8Џ�
�(T��,�6��ε*W�3�����.���vC�A%Wy�$����h�O*ci�k{�e����U�=�G���!ʺZ���ir#}���0(Y�|}ͩ��C�d��z�aB�c>D#'_����&8 `�V� ����ma_���=�����&y/�֋�0`i�rC[��MQkP��D�M�*(6����퍖�x]c\���hZm�7W�V�����ܨU��ሆ�9E�͗����0d=�0�#{t�iՒ361�)(��N�MQ����3�p�Wx6���D��u/�����ho�2���h�)"ۃ3����2�����=*s�<�H��N�1�Xt�p0�NG�^D2h~�gg��F#���p::�e`cơ	5�7��K� ����KQ�P줙�/ 1K���VQ��a��<����V$�Ti*�?0�2'�<�3�3�*�J�e�q�ʱ�o�Q�R�nħ�������٤!h�ʚ����� ���>[|�i���Y)�:�Q);�,��xr�<B�#�2Ţ��"
 �_iȨS�jv��2Y�S��X�0 �q��VYĲL�()�ظ� ���T�$�G�vTuQ;���f�G����ᒅZ�''E~ҹ���*����Ɋ���%�I-�Gՙ,
T�h���E�"����� Ёp,p#�����B��NT@�'hn	 ���-XC퉄�K�)��Z�<�I}�QeJ��.AgI�j�5�o�|&�t�d>Q�eȡ"�ʾ�J�4�é������0�1pI��������e*��W N���S�X��h.���GGfV>��owy�!f�
����o�pA4oѢU��H��nGǑ��g@Br�/Wqf��gQ] :dq��=M��Iisy��2�^<'Wa�'�/)��T7����?>.��㪹 4��,�?��=s���A���܋���L�P�P����J�vc	���GQr�8���p�dII���"9spMdo�!*D�".�|�]=�⎧����kD�	�8�3���ޛ���׺W�EE��\xG�6􄬑j�*l�q���������B�Gw���fgf��	�5��ؕ�k�P���YEI2�ͻ:9���;���xsG����N�z�NZZ�e���s:�#S�}���Y٣o����IS�i��7\6!���҇�y�I�$Y��ѐ�AT�pc��!M�Un��<z��i{�u�t��B��q:��^�=�a�Ӥt��=v���ћ��)0'ܪ�5mߚ�\���=�2��r�NhX������r�D֪z�x�H\�Jw��_S��{����U	��/�)"c}���>�,p�� ��M	u]�0֐c,�� ��<�����",�S�r�Z�{���8D����h�\��ܫ�5��c���Θ����1%�i�6�&�r�5���7����ks���X�t!�߫�B��=ԅS1�-z�n;Fs���W�)b����Xс3v�=���o�P��]����{+k�ߪ�2��l����^���:���;�^���]v�o�����f>��"2�S��)�����9��
�|�,������xzH$��(�b_��PƧ�y��g��X[aWN�-���f�hlW;@�%Oq0�B��(N�X[u�̜�o�2m�kg�zǡ�]f�f�1�L�s
^�hiZ*�[l}3M�N�皔~n������2�FLz�Ǻɭ/��K4�*B ����D�5R��ﴧ��2S&I�{A���ő�E�#��9�jƦm����z��P~�N,O8�ݸR*�h��1�� �b�2�`*ݝ���'x9a�YI�-��s��R�,\&�� iV) Ea��˟����'I�6�r�5.�^��mA�@Ĥx��wdK�Ev���.QK�T���_��:Է|5G9z�"*�j~�B�Y��چ�,H_۵�2�	z���`���4W��?�X%�������ޏfvh�E-s��#��%v4z�up�,���ZJ�]���ƯCN���m�Ɵ�˓V�z�rT��y9�e���5�;C����ЯS�^�S�k��P�V�2����i��ҿ�b��l�z���gq2)��4�I�������Gz����E�L"2G��\K�Z��⹍ |��秌_l��|��[�j�|�>^Č��l�ڋ�,�Zo[�[�@2�/)�