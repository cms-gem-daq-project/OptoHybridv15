XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o�g�ҥ4Ƭ�!-�����a��H�A�ɜ��5�ʌ����_g�t|��"ܡǱ�Gk�
���x$d��_���e!eԏ&�w-�[~n�WUL.;�� ��8c�y.\�����ߘ��.��S,9�X��{dͼ�l��)�5����JV64n)��n~�	�~�MGo��]-*4\2d�~f6�?Q��"�{�\��C=��%��m�n��po�B⧣� ��d���aW��E5c|C�8A�]�� �4�*aޢ_;�n MV���� v��e�4�p�T i�N�_�w�9��[�G��i��_�t����6>W%Q�
F��*��U�C�r*M��j�x%���Fsy\e�J�a��ʜ���pUf�w��"����W���k���v��M;�ܤ�_}Uj�pA1�&#i�Oo
_��%�8�:^�{\����;�9��f��$��Y��h�j�3��ఢ��dT	��w�jg|h��9��<fG|~"^W$�' �}r ��'���h.=�����sÍ#= �@�r�d}��������pZ��o��-x/`8�@,,d0l�d����}Jp����;a�A"�!�wV��EL�b2�%�7���G
F_닠�.�;�%ƙ��s�d�>��H>��p.�Ǐ��������������mr��@ђ�8P�h�s����t�Ut��1�_�2NT��{->�$
ua�gc�۲Ht߃�z�d�R�m����K�߷�!��Z���C18����	]#3kH@8W����!'N��XlxVHYEB    4a98     e80%��f��n�ʹ����"��JDT<���n���(A��6@&?�ps�:��P����8P��3��0�g�ls�ُ`��v)�ͼ�&{w�O�|��yR��{���t�z�]��Є)FS���k`��¶����B�S����*��m�&ܭ ^g�
L�JL�H������x���me��vF4ܔ3�p��~���NT���z��$8f=^�ʐ��T}���k
�QIv�(R��S�JH%0�U/	OSH���-������/�@̕D{�PTV����.�*k�z�s�|�
�5�2 O�����A*�"�C	�%����f�'���n��`<를k�]2v�I���ً�����h��R��]���?$)����i�s��6`c�ڢf�Z7����q��S.P�|�"棜���DܳI->OQ����]+���-(u��7k���3	9��)��?t������%�4�/#3�������m�{ySW�!�6�6�=�Z������ԣ2���`�'5�D�LG��9v�>�kA>܀���$�
 T�0���vw���>lWv�6"/�NVQc�����
��V�E̩����֚���4Oxmm��^Wo�ߜa�8� ���]j�Hv�%:<�c躋��<�%��Pm��`�|��}��9o��x�;짺&��S��� l���&�V��H*k\(��m�מ(��pޣ[&��ݭw�@��mؘF�2[T$~c�Vj�>����J����E����i�M�~���T��D�bW��+��ذ���f���m9���ᕭ�W�HH��o.n�p� f��8�fA$*��pn0�@ ~�٧>Ι��k.����0���V�hLvZ��¸T*�^:���ܯ%����#��0�'Tʏ�)1���'џ�aoA�&�N��S5���?x?�=� �&��������A>��Jk��+���D$�߾�ǡ�Z?��r���_P2UtsF���/
�0bW&j��g�El������h�	{Ƥ����ʇ���zV��Ւ�:I�$Y�\����K�X��ކ�zkpq��+�a�M�(�r٤V���P���F��#����Cu��ZB&E]��t�"�b�B��¿kd�?~4K�9��V�1#>��M�út�؊.��4U��s}e��73U�C��D��.j�u�¦ ��)�YԘ��/o��|�U�K�'�G�m��l8�ӟ����Ɍɍ�4��Ҫ	��[��>@棿��S`��O��Dܕ%)8?��+&��Ld��I���A�,� ���i��i�D�@�9l�wGb��-S�����A�\S�)n�M^��0Ul �HZ�.�p�����`�:�������
�.���U/{���I�q��-[������h�AB��0���	��,"����7��B�}$�|��*�)����IjV�����I�j~qg4���+�̇��-�I�7���K�{����B����(~�:��g
��t�8Yx��~��B��PW�y�q�jW��1gĸ�����_q<��z��O��(W����B�����CU�e�
�������tR~��sj=X��#M����{��_����;qhkw#��a&���5q��Ә�h�ӫVMp��}��6��D#�#1�~j��}Gs����T�G��;�����?�R�FkL�󩳩��jl5��
�u���d��1[��ª�9��W.�BO��Q�[B@1��-s:���Y}����j�Sk�?٥���%���tp8T��u��t�2�����5/B>��2U�=�� �����&�S�6p,�BH���4|���β��ֈ�c���M� �ݽQ�kn_T�LDڿ8��ձ[A��#:��a���X��叾����n��|�����V�|�FIĠ9U(^2�\L�`$l��yk���Z�,�ӈ\�?F��^�o|�%֦��r��zg������X:!�Od��zvō��	3�`�0�X�'B?E��I"������κD��2���J���Z2^� ��/�k�PV�P6댚5&��?��P���	���v�-j
�]�fK���#�S��ܖ�#��k�0��.�����0���n�>=���K��ٹ��T��Or�O%g��n��9��b�;w��7)cS��K60��K5s� x����|�ؒq'w��ٗ�>XSC�W�)cW*���+t	�jQ����6Ӭq���~���y
����*�\R�bK���I<�tzy���$�c�݅;�	��IJ��Z��=O\A��^hw%�]C{����=� &�KxԳѻ�������Q!����⠯�=��	�"_��~��?���/�z7��%�B�E���Z�p[�b.����}D` �r�|[5hxO�w׭6��ȳ�D^�`:� �Ԙ�p�[��6i�tw�٭����'ɸȕ���A���R6j�s���J��e�
*��x����b}	#�;�xW�-����k�_v��pEţ礸���T�N;�Di�m�n��`Sqy�'bg<��8I �n�b-���U���x�#�;H^U>��[E]��'AU����n>I�c��&xh��3ߘT����� �z��f>���c} �ݰY`�m���cH�މ�v��	��\V��������J��䝸�{PN���oa��Ril/M�=]���W�?�l#�d/�5�D[	��`���F�-	�4���+�%��0�4�8ħ����|f�>�*iٳcӁ�^O�%��������=ٺ�����AD��xvIJ{������˫��� �2�u{=��79��#Q�����H��z�%ث�H��$�����3�. ��
zKj�����i]��;ہ�v6(=�k	1x����T��m�ߚ���.%���Q#h�w�je�nYѷ���wR��|��!"V���]����a��?҂)N&Hut�m���HI )Ļ%���)��~��4��B��,dY��>���3T���>eZ~,��VE�"`՘�h�lĸ�:�o"�%�c{�'"���=u�Hv���1��φmp�\�;4���/�^H��p��o6I���m�9���b��Ld,�D���7�"1�q�P��_����"�z����c	�������l��Qzex
G���^:dxL�G�����5Mp����W��]wLz���g$�:�1����d��*��*j�B ��p68U��B/暩
���pd'�fs�,�EѰ�Z���s��#�؅���~8vғ�9f�܏�U؁���jq n|�5(&y�(�^�D�� ��e�����K�.���B ,c?�e�3Y��A=�m]=�u8܍�����#20��YU�6"�:
������@D���iM=��a 3��~ �↵�(h�ч|gy�xp�dHr?�QyCh�-2�������t49�i�TuТw`τA��DV�|��Q6/�Z��⪢)dB]��Y~H�"󞿓����"SZVgCD[A@G�l�R�o�-yc��-rS|C]�ӰV2��C��!�����O�ׁ�Pz��AZ�ε��>�t�F�s#7n��W����S~^��"�AI�qpN��q/(qe�~!lyqS���DX*�u)���4d����;��_��
坑���0}Z�3B��|jƕ}P1}Wu^r��F^�q?��{N�:>�iJ}�%=4��v��J?�4�i�H�{�