XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���bq��C
�<�Z����{��%e�KE�7�V�n���ۢI���o�&S�%�k�y�K�LH���I��K�h�);G]H��QX�y��F=�;댹��B�*P�0AZpM<0ᾐ����NS\rߪ(�_e<��#��m��"����񊨹����M����U��][�W�V��2�Hq���/�7Z�����Re X���~�WDN�P}l��ij�l�+�j���T�9�a��0�D!̶(O,1Q�Kuؕ_�1�0˰?Y+�n)���B�U�)4��˂����w~k��U>� u�Ր�A�fϭb=E�`:��VfdC�0g5��H�Oޕtc��:2y+����ձ�h��I/jAX\M��i���B��quJ���!�g�����c�_�"Hӂ�݉�9�g��H��.~��mR����gc�>%�o���ʜv��8�|B��p���(�:I����wH�+oI�
w���)�æL"�4ه
yiSƛ�˰ �_ʍ	��g�����ܯ7V�v�T�R<����w�cq����Q�wH#B��ħ+�v�e���i�(�#7�����^�4��sb	�����f��ЀtW�v���h���-T����p� n�<x���V|w1�/&e`]}�p���m�wU��Tw�9�R��O��� *m,t�!>��cڬ�$K�4P쪎	`�.OR~�&�4���s+)38��1����$��b�p�����&/�?�2��6y����V�'�=�ԕƄuYH/xV�OXlxVHYEB    458d     8b0��n5��Č����g/<������'mX����1����ެ�pqL(1=DE�gs\-�%S�L��7Mh�rt���-�?�0���[]�CTk=��nT���k��U��u �K"N��ة �`/Jڤ�V�%���GZr<�ɂ�� 7��2�Ic�hЖ��5B�����̻��1u}���Å�H���� 9�*��Q��6�����t�%f��M�"t�?p�u��B���z��/>A��������-J�p��م$!�I$��s��+��d)3(�g'$�t^�XK�J�߿:�+j8G�8^�I��Ue� .�T6Z�\s~�F�X^sǛ�4�v�F�r��q��i�O�м�k���sLK
M'�]M|N��n��u���3]���ph��YV�)Ag���>��>佃��2��^)�.��%��s�7ͨ��#Cθ`Eǫ)8ق��\��'�r 4py/���!9"���SOy믩�%q���Cy�1\����%�:��C�4Tjk�b�2�n/��L9����7��i+O�Ϫ�H�>���M03�q���8��>a����6�y�ɿ%м4k��πXd��m0�Vy��yt������$[F����5Z_�1���Qn��>~ۏ�:�������d����Օ���t��p�]6m�y�Ne(_��
��15G�#��ɞ�L}�`s7�p�^"{� �O���,�6�Y�3k�M�b{)�M�����`#fWl1�_�¹�2~�>�R�,><D�)~��U��:V���T�50�F�O�i���p�TK0Ѯ��l>k+*���Ӹ#�[E<��ȭ��N�?>_&v��C��j{h+(���2�x]��5'+v���c�Z�y�ȣ��z�2�q3\����E�D�*�*K~ؓy�p(���"�c	�"� ��:���8S�9�9�~��8a�l)�<�bɚ�����}��pم̹*U�
SJ}NC����	�9~����s|K�L_.d3~X��ı�h�+s�M�|\���aǐ�6&�e+k�8q�k�75��H�:4w�y�4C���u{=*x���s'��l�TM�1P�e��&������0��f�}��8�����Ey�!+�����$����6� P�#?݈�<+���U��;@ܻ��ri#�Bn�X�/���#���׶�T�1-�W�.m֦8�U���7��ͫE�^7���+(�7�|ϴ�F4�\�������J��j����?��I��'�ܰ�d�j\b,e�לEea�l��=�����J�������G=?�����
#��8L[���U�;�`�I
Q,cˍ��['+g_J����I��Bo�}SM�$z�pC��Z�x��]�̓�7w�6?�Y��I��21:���Ɯ�x�Ž��v��NچK��*���O�wրH�ˮK^LwXhӊW$.����'C�-���#��t���TP�m"��H�mI��6�`+Y�,�
f���Ͻz���O����c�[qo�j\�Z-�>����lʍ��Ye�O�����=]��F�l��v�GZ�)���%��ۄ��S%������f�(y��hE3��1�~�ڪ�8�;m��fԆd����C��\�,j�9L�)��`0�u��J�i>k���C.U^�^��'�]w�p5X�ā�>c�d�yNqM]ˇf>���J��� �k#Dъ��Z��4�_�/�-��t�;�p-����F�YS��������?b�}Ǉ �§��d��`����6%k��p`qJ�վgG)��W�	�CIڞ��IO	�-Dz������K_���eU�s��p	,?�j��Pe�T;�2�ƴ@8:��o���1X֫V���Wn����e��ly�,��]"<�y�sS�a�7�6����g��=��P�kW�:徘~*>�%��1��2��^/��t�`���r��W�/<-gޭ`o�FW�1l-��d�j����������N˕(�LQI�BC
ņZc��M�=���ıL���Ȯ��)%('VHe&�U�6�l�T��ថv'G�������"M�vg}L)�����	>!�/{L[Hu��
}�lC+�JU,]*�����I��a
�?ʺ�^�4��u�F�xĊ�D��&���ݜ�Ƨ:�=m`n�����X>�*/\9_���C�O���%G~YH�h�"�5�s�9�Z�L�Җ�]�y��&<`���: