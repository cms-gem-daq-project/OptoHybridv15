XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�s=�.&�u���I�Fv̮Tc'��U@�r��R�|Q��b������$��Q�6y��IMQ��~����M��ބ�잚D�s]����O����*F���:܇�d���ʳӺ���v�8��(���e�\�8� �˵^��U��Sb�E=<�ǎ�4[)�����Z�H��VP�S��ʟ�	[n�M`"��r��C(N>�L3�wV�.�����5WQb!i��#IlU�KHLP���T��22�w�z�Dڜ�EҬ\t+"����,����{�$6�k�M��+[��;d�P�O�h�f?�J�%�!B����M:����o��Z=��鎒��MD��&��:����b�x��c���{�A�s�
R�$�����ߩ�F%���X�2��1ov�/�?9"���2M�;.�����չO� u����ߞѝ�IJ褡>H�-㌏5:���1hg�?]g�K�?2�f�Yovp�s�g+K�E:��RC:8L�_�՜��Wԇ~���t�@�+j�ᯐ�(V���U`�O
⁸�<�(:�M��*�ֆ�^��ȳ���2�<N_ l���ۼ.R"�����&J����ܷ��l�8��<�i����uN�м����Y�����)"�%�t�J��Hu�a���7�2�I�`��/���������<��t	���Dl0���sd~])s{*;�������L���R��9tS�G��n$\D��$��%nT�1�0��"����F��N� �!�H���7ayXlxVHYEB    2816     5e0�� W����q�d�[���ٯ��vYrS��j�66��M�CF��G�f��0:VuA�����s���f���B�����@�!���Z@a���O�� �� �F@�+LQA��b���S1�%.ˡ3���f����hr�9X���p�t��V�6��p�n���M`��P�;S��J�qZ%)��l�Sn�0͏�n�F��G������@0	y��q}a��L#Z�I���C�^U9&}�p���p�OkL�-��)����v�����'��R�8�̅�n�"�5����Kb���*��]����fo�`�F�W�aAr�JÚ58��&\�	�EX����7>�l�q}⃛E�x�2@T�eT��Ƀ>���*s��yN�~	GY�͒��r^���(���AU�0�"�!H9�z�����K��\����'n,�e_?ܚ�?����*��M ���bU�2nç)NC�c��ٳCq��l�%�BZ�"&]�����#���>]����p�q���U�� � ��;2��nD�x���{���\��~�'����H���:���:P54������`�_X(���^��>]I��q�ŕĘo��;]�`�00�r��ӭ�e`�V�]Sg�]�@�N&�0g�Ӻ������N����=�櫲�/ƍ�"���޳�e{;?v#�Z,�P�HgQܓ���&��5�s������^t�^fgr��},��ڬ!��ם���WX�]:EZ�j6:�e�eE��F��14O= �q^]F���V�#<�ر�~�O��:���|���&(�)�Cfx�1$�0�d���nx�@���t/��	�x	�E��
E�L�����)¸��w���4!1|ߡz��#=0�r	�y�u�w������n]NΤKΚ#����z���P��/��v�x-F�F@w_Z7�ev�N��:���5�\�9�AŔ�Wo� 4�ۯ
����_݉;�|��z�`N蚹��˒������ }
�q�ſ��m�ᇜ�JbCy�"�gA5��qh�DEB(��{��{�ۥ0t�Ԙ\E�0��?r���0J�6w�0��aEO��<�'wz`+�Y6�B��i�;Ķ��礗�xA������
V��禊%)�i��0��}�h2W�|F���W�G���W�()&�N���cV�L;�_=����%��[)h/^;�T�rP�	R�|�竝�u,�f�_�"���o��t�?!N#�tD!���$�y�z�^��)�1�-��;����[��8����}�J�����+�?���gS:�+�,s�Q�u{�מ(H�y���<Ʃ�`�7w|<��hd��G����~�Tg��0��� ���N��қ��Xj���!r��-��`�N�P�R���\^\��0��S{�|��Rn�=�lV����,��rY/-k�|r�ð�|G�DV4W�W]��c��kK�3�
�\�t�؄�|�;�C�YA����!r1]������q���r_�Ax�N��