XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w���ɳ��Հ������u+[������}��r_�A� CZ���!k�R
5faD!泖�߭I�f,a>n�ò?R\�91�b�!>��{h�U�3�~����*��8"��+~ňt��)�?č�0Ei��C��
��kt/�uu�z�3�v{�p�o��{�]���m$���� �6fF��Yz[�s$�S"ΓlNÛ�3\���E�@�$��Q�`�)��:AX�T)�3��=�;���������:�Yd�uZ�:��u�&��.4��Df�1�0����q�V��ޭ�+N�T3�`U�ҧ�	�O^���(�t�ށuv �f�SI�)YX�$���� �S�Tc�[k}����&GYHhy���!���q����·	����>��g�4��I�r�A�v��E-_8�̒�AitJ;�=TB�B"T�P�e;��}��J ���N��v�������{��.�3��aV�p�6;]��>�p�I����}���K�G������-u��'X�<���Q��a��	
up�n��'~��iҰ��(��G�1��6F��0�%]��I�, v>��,����Ij��a���1��j�W��R�ƞο��_�J��;��Rm �T����ִq�?޷_N1GL���7h������� q�փ��3��>o����9���Ns�a'.��a��*��,�5byъ���S�$���p�>h�Y�P��1�1 ��W��7�;w��r��K�XlxVHYEB    2d5f     800=9yP�=�;+�8Y�A�-�&8�9す�w����[&�����s����7.�v �ҠjbR�ڭ�+r��O~w�����y@I���R�n3��HW))��Z6�F��֓Tη��oK|���Y�Ay��Y �>j��a���
�`�r��<�n�r���5�v|���ǭ�d�}�!7�%P��D���e����y��h2�!�@MpB�H�@�WK��X���0l�F���U��^��KT�rB����tV��x��Y�'ׇ���'u+�k��"����$k���Pe]�2:�S	��|��TV��i{����g��Z�i�|�/<��'��NvOZUz�����-���G?nt����/���������a�����H�ux��T�:[�L���3�R+s��n^~!�|��x���@<���܎Q	ܹ0�<D|�o����A��6�˿s� u���G�Ԯ��1r}O���ė(���\%ͤ�-,���*�����5�,C������<$��^�ke>�j�S�m�.��~y[��S!��7� ���ã򎦦 �.L>�}��%�e̊�x03t���Sj'%��]�����2������Bbt�<lϲ�/��h�t��\����O����ޣ�\Ű�]����hfg�
��� f, F&�1�K��^�M�O�-([1�����:��x��	ƙA2=�%�P��aZS��XU��@������Ǥ�ZT�t�FE3=0��HcT����<β� ���d�&��:t��|�����Z!����p��yǆ|�}��=��?OP�nЕ_��-	7���R�����Ba<}|0m��g@�e��"�E����l��S���nz��d����ly?�j��C��W8Ew�?�K����^�.�,H���H�S�\�I�S)C.,�d�a� ��^KN<�CVӦT1�5�YM�\�C���᱙��Ҡ��܋P��3�Cu��S��Խ��h ��B�`~�[��
��#S�>���z;�/R�^C���[jH���><+ߧ}B��$�U�*y��C���4eZ��n
��h��?î�0����y=�F�+�kz��*���ᑎ��-@�/F�s�V�g��+@��E/jm4�������`5XRv�іR��ď� і�w�2�P��0��Jr.��|{������D�����Łi��gL�[���ӑUn~%%Ŷӓ��2�\�{O���JJ�w}����TA]i�_3��B7jT�������d���G�74����I�5@ܗ<��e�L2����j�dZ���|�pjY��9������\�,L�=����G1��K�1�WGQMTxꊺ�D�j%��-%�Ϫ��`��fHo�~�-���fJ����:W��wc
��@vߡÎR�8��{"z�4���r%����i�֠2�6@6D��Zy?X݇@�.����9/��aW���֠%%M�1�����)�L��x ����e'b)E�сxA�@��{�s�����	v%^�OV����w����(
fQ�V8��Jɺ���ܔ�kA�H�*����f�@$I����GҒ���y�ۨ0��ce3� 9�H>�yK�b?�[�6$c���pȷq�b����Ͱ�39�{�y;˞�W��m���Cʴ��Ǫ�xV8�c>����<uS$BV/��;&�r9�� ��W"E;f*w��ʛw^�)0l���e7�/N��a���_Y��t�H(,��������{�ך�7��G(���ៜ��}�e�o&��7�z�0��X#�Sp�]U��ۿ����u����9}	ԶL�v�R��\��O�X�7��6'�3@/���Zߴ#Nh�����&�*�*��g��QX!}}ҫ��$��4�{ސX�~|���'C���Нk4泮��i�;�ޛ8��XCe�L�-'��{R+</]��NZgמ�}.��k;]v����!��ș��B�L������U�mt����R��+�T��.iv���8PV9L�Z��;���