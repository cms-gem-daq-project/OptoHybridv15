XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9i�/�,�>���r��DU�	�E�H�$9�N�d+�~'�A�� P�y^��k� d�m�a'bB�<\W��@��T����a��k��n���"o�zܖV���%�͠�������$@\��}U͙����aU�kV��o�!`�8�<r�?C�?��r6Wde���ռ��g�.��I�2A�V0���~�՘g�P@�)��G�kl�wk��?	&���{ú�Q��,9�۪̈́�(&k���K�XJj�a�ds%w֎2X�$���Q��v�(����d���Ц9��ў��� ��Tw$5�n�>����-�r�=|.��#Y�\
8��CS}�٪'�ì�7��@ ��Rfʮ�.����#l�k|]� ̷o���(~�+�DY�uc���{���R� �r��rb�XES��L�ҏ��[7Z�lV���?�uh)����*�����e��ٗ�s����b�K6��=�m�t�8T(ޮװfV���J"�PMl�Ք.���x=�"�{��Yܭ�zf|�����M�ӂop{�'����-l;/���z�p$1��&&c�kŷ�da�$,ϯ�+6�Q�=t�k�Wv�b@0�CV�2��U�x�?q���ڝ��)�Im:���،�����eh��N�N��y3�h��鴈��X��bW�Z]�z'cPӧ����K �I��J�P��=~B��C�̀P�: 	t�P��r�[�ojj������µ��o�}U�Ґ�~z-����*"�5T-ei�����XlxVHYEB    4b0c     d60��)�ea�a���jYD�;�^�\�'�/th�^�ȹn]8�_���j�gz��cLw5� Nu�s^4ǝ�����w�d�����$ �W�:���n`�|:Y�{���	v���N!�ɫX<w(3�>����Y����t�N��4���L-���+�bG.{������t}|��b\p�$y �x�nAz)N���Xͷ	�h&������b�B�bY3Mc�wlʙu���uy��hL[I�^.�?{��y�
�K:>-L�����;�s�m����v�e�!!��q$O'C,7F�|ً��&-�$|(�âNqe^����1�%4�<�hQ�m5k��0�1��������K\�XW<��X����Ɗ��Ʊ���}�=�R6$�Y�|/J̬����d�2�N"�!U��	?̀k�9�4IY�
�t�U(S��f�U_H��A7sJ3��@Y�M���4�\{�2��W����އJ.C����ɔu�F�����O�Q�?�����CY󑝻����cÊ	MJ��2�F�0>��t�)J��xn��!���(YX��0Sĕ��m�ܲFJ��K���;�IX����\!�(ъD���x �1���-��H���6����]G�����)kf �gX��ԛv�o�D��������KH@�����q$�ۊu�=�˄r,�Q�đh��#N����p���	��^�N`,l�]��v���RZ���m$��j�ϯt�	څkA�������:�C���d�h�n q�<YU�H9�?�/ߜ��!a�S�m�*1*���(�N�-݆�t�Jz@?o5�8��rf���b}�s�����f�MU{��Z5i�Si�]N�]�O��i%K�����u߻��>�r�`��|�֊w��b~d�eN#���j��Wb���(���Q?:iWy�QFvS�	���4���8�V'��#���Ө����%�/`�[�RO��J�����>Ͻ�_��OE�#�wRD=RA���N�ڡ�9͜o�DOّ]��ҽ�>�]�T�n�Εn��.v~���,������-g-�R��y��͙�K͍,9V����cp��(�u����5P0j�"�5oo7�y��[(�jth;%Nd��� �i�1�jk���5�@�l������I��y>�l?؉[1Y�s?=��@��O88�x1rTb݈d
�@[�ݍ�O���jw� ��gjL_��L���
��/P�/��Ȫ�<ZS$W�ٚ�������A]��;��sg�psgGy0}����+��́V0c'��{V��a:庢�šn�������bG8�X�����,�?w��Az o�w*@�ܜ�r�Xwc�8������N�
}8�I���W�s���}\�M���ش���!�����͝f`���)��'����-��yQ����ŦV�L�}9=���㛑�O����8YL
��s����S����IIM�R�Zc�7�F�`����~�=P�z9�rE�9�!��X�YC��.���T�I��=�M��wM����y.��Ĥ�3��u�T �@W��AEj��B8|S& H�� ��v�I��P��#�p�a�~��lJuYW��u�a�^PnZ�^ ���![ #�z7P��Y�R2����Ҡ@�_83��,۳�dA9�]�x��~,uA�Sl܀�h�8�-Fd��Xu������o�8���1�F���(�iE.y�2��=�X�NK/��;�L�9�u�᪑*�!��'�G�M��_�d��֌��Kx���zg�
�����a�bAm�	��?���㣐3���f��2�j�VpOm�
Y� S\��Ж.��@wSQ�l��5�V{g?[�����BQjt@�]���|&^�·�'cܥQ���\@��3����o{����I��S��Hp�&�D��]�N�3��&����{�	�N�F�#����:hs�W��K�6���P>�n��¹�����_����g�i��w]�D?�o�ޥ������	5�9�
�:��k��s����"���B��r��ú������bSL+���ނ�#"���i����6ɰyo��G���Hv����F�sx�buY�R�V{:k,�8��h�Z��}ȺǨ4�y��=*6u����	S>L��1W��|�����y?���u�F/�4��HТ�R0�ZA��p�+:0\���M���/�t�謴�>��ۦe��(eOE툖�(��ġaΐ�\�V��t���nТ�dШũ+�`�S��6ƺ' M���~FETc��F�F��иc�"[��7z�(��u|	�o�^LbJ����iT_��c��j:�+3���?N7��`o��S	�{%vA�k�ם��ܝ�j��&K��'�0����̸��{N����o�%��X-\�`18�5�T%�b�;Wd��������t]��1�u'qa����7� su%^��@���yޮ6��o'�=����<�.m�m��|�@d���L
������J��S�m�O�15�2�`T��&�A�`�O���lrgF^ �?Z�:�
cI�|jc�W�wZR����/��U4"�by�7��j�#��x�'�A-����Y�Ȥa�q�C`�.\*�'�M6���?���
�oF�����-��d��	�4��DF�\��U^��$eW��ٷkz�7Pwg(��b�
��;�JD���O�s��%r�v/�v���p�Ӿ�"~f*�����Q+l�$���n��D%��*�^tXl� |᮪/�Z/���e�Q�"0)5A� r�(�a=�>�%��/������#�Hm}<���@�*����-J��xd~�DE(.�F��]ˉ5�	p{M}v�z�:{Э���o�=WY�������y����q�	tgۿ�!I|�"��)���	�^��qz��cΕH�q�)%b�/O�"�vr�������%��>8��U҆��Rm<S�_G^@s������r*䞖Q���'�ɝ���]�>�Z��_SL�	a��zD} ����Ax=�+Y�D*��IP䟑/��O��T�F��<8ey�9�끛=�F����ӥ�Nx?ex�j�7��g�[��Q�x�f�����W���1�5ߣ��������b�t�0RT/��O� $����n�h��zKP�m-���6��Y�&9mC��/� ���� v�xp�Aq��+Y�07��_��[,P��5
�#\�+`K�azmy�C�ҝ��V�E��u���×}��#ɉЁP�E�ھ�v+[�b0�i�ZY�-7��tK/�o��Ns�{^�ݬ�ْ!����]oz�K��ǔ-s���ϊ8��[I)3�A�c?l���y����O}�ĸW�	ͺ� ]xF����������L��zۤ����}�;���z����E6y�h=cn�R�W
q��