XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4�"+��T]~i�H�&1�l����Y�����]��P���w�s�{�y�6/��JrUV�L���{�3��I�b�x�I|�#{p:�B�`nwً�E���J�Zi��mFu�Hhi��'�xz`�xd�Q//�Zǎ�G`����U����=Gi��E��k���P��u��9�ק�S�>O|Q��f���M1͔.~8}�iNN�zH�)��!�(&��s��K]��0���.p9�w5��9D �Z���]ϵ7`�b�/��q��X$c���L��+�'s��9�R����TȻ��Ʒ軿w�bx���cD輦����22i�z��;I�"?���9�����CB��))��u��mS)�����b�m��:��D�Ǐm�}`��,` -�a�ϯ2&����M�����A8��v�z�\���W��{)O�"�w�'E�v�� �	�-c���l4�����P����|� ��&�R���6FF}o��1���*e|ݼ�,
݇YF���5������^��.���؝��@�_���m# |�����_�.���o4*��5e���Hi��gծ0�$L�͚7(����,��������ޤ�"D]��CB�ǚ�nF��Z`�R%�!;��L����Ec
�����$<}W��-д��y�+��h"<��vЇ��2r�C�Jfo��g�Γ�[й�y	��W�|�d]�c�1+&�M>�"=����x�k��W��`�<����H��c�#�vA�/��L���XlxVHYEB    152e     580�,���G;�Uad�J��s\�e\��G�l܋�V�z��V��-K�HV�s)��\�s�(I.?Sa� ������x.+�/O> ��M��RL�-�D��Cl;.E�Q��ɰ�R�P��"��Ia^Z��}���V�Ŝ�֙�#-�[jt��k@X4�!�qwL�qX�˺3�*�-�?� M��$˿��ʛd�~���Y�uToc�S�)a�a.�L�u�l�	�+
�RE?���KU\d�Z��d��9Ǿ�ZW�&1z�ʂG�<����3�{MT��-^g�Yi�]�=;�<a�Ng��]%\�沲e��7{+���![f�/�#`'#��?خ��DL�[�iV� �xg[��Ը�]|Xn�Ȑ"O�z��n/��ӆT6T$/��R�b�Hŵ��Cyg�0/2~�<%KցC�kj4��KD��@��m֓m��Ma�+�p0I����2��0�.�8~,����( �\����6��5�0������.@s�LT�K��ߺ
?{wr\�B��p��^��A� <���r�u�����v,�b7Y�n��k�u����]���쇖|xP��ڲq��&kh�Z���_7�l̬t�GkL)CU �\�)�/Y�cW3=��>z�����#r��h��L��VW�v�i���*����f����J�M�lj�AU%�/����Ô.�8�J�y�z3���%J�����`(WJ�t��V������G����k8^(}V����I\�C!��������n7�]�H��8a��d��[s��\�z\=c���.O9�"�b�=y--�>�G��e3K����82�lΓ]���}���'�F9 �_��|��WF�xA�<	���ӱ��V�H�����5��'�z�SȚ����2���6�qi��g.�E�@�'h_ோ{}�����
aw_�^j<_I��RB���
�O�2����
U���U		��,��h]�42��޷��s�b~j	yʀio��&��sN"pC�޺cE4�7kKki�	���F �̕��K�*?_��軔��#b�nXd�ɿ
ծ���Rq��H��7#)��x��������Sy��Mn�"]�{Nf�C�g8����q������T1�d��jq%�s�\��E��s֢�����:4*W<=n�?��E��s�O�M0b@|���D�y��%ۧC����,�"�0$�������N����VӖ�����j	���"q�r�:��F'����Y�ƌ��C�ʷ۵*[�25�k
B�q%8���`GG�Ӹ���b���J-�h5�����A�b�4�� >e|�(oI�zq��9fr�P�0�s���;�+�vm=���G4��n��F<a_����j@��e@�