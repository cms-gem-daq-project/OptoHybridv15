XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|������k!�^Y&«��A-�P���='��1�3����v�����Dߕ�㜤zH�6ʿm�j�~j���O(���:W��/!�u�ݞGD�k��+����4f�hI�(f��1��-0NH̘Gr,:�"�y?�bS1����\��H���g�3�P�p��������Ъ�Q�4�b�&�k�'o[��q+�����Qd)G*: B�:3�]�D����`m�9�@�F��z���ot�a8�D�\����5�z�: r������2H����gٽf['\�ig���\	蒷�#��6A`O?��7����1JUC�Z񸻁<�j�	���a�7�/T�)�K�(������f�������x��n�����E��%���Zm �C�1��&r��;���_�@!����I��v�8�+�&���z"W�&�4#|�,C*���>��Ӭ���0�S��E�f�k���0_����N��x�N��5�4��q�ӛ)]���&���JZg���	���{�+)�x�	zY�/.H�;嵉����$O�9����H���s&L��eA &����ò�!���E����V�;�^��1>�aђ'dۿ#Fn ��\�B˄�_s��Ir�W|����@,�S���{��wb�lYơ�ЎYŨ~�6J�2>�Wۥ���~���I�x����"�"��{�~J�Uʩ��85�1,{���WBnU		�HfV��M=�L0dh��7���#�h�`4���^J{`��XlxVHYEB    282d     8f0�2�������6P�>��Z��e���ؖ�p��ٿA"�	o�=x��ȸ�x*�� B�qf�����f���p>C������@��7���!�Mh�����q�-���V�
�M���6󏚉��z��h�$E�8`����M��M}�Xm��i\s�W�y�.��n�,ȯ�n[���#�JC�|c���.
0O�RG��r|U�<�V=��"�/�E4��\htRB�w�d���� $=N�Bs���#�4����Q�+��H���b�i:�1��c��J�t!���se���Vƛ~���}�Ͽ/xV�ղ�ʀ��T�V7J0���C�B6M�r~L��ܢE+� ���O�[ c�e9��s�~%�����#��\d����

t�*��`I�E\�:��D�����1����`��;���y �����x�c�*�9~���-����f�x�m��66���U�k��%���~*��r½��Ka�iH�0O9��,��P��x�7�q��Pe֪���Y	�w�꜀'���<>����J��A' �	z�u�_ް�)�vC\B���i%�^	8����9'� a�.�|aHWh��>��F�m1% �����Q�c��V]�c��uCD2�VX�}T8��m?�3K��?-b�N�m�%)OM֊��E/�D��wz�I�׈h�&�:�7�q�L�ɴ\Ǩe��*��z�m>])�M���mUz�=�yU]wl冏;���(z�_���#^$��!����1N�tk��og��88±Lɉ�<X�����S���Ew�+a[���!�!�<�csx����Ɖիzbu�~�p\�<����d��Z��:����I3��a��� p�K5斑nQV1�b��J�q���"��F4�����DHf��]���%РhG��?Ch�[�@����b���V���ˠ�pV�ˏaQ����@Q�_7Q!$תΎ[8��?S��׶�@D�6��ԛ)<C��₊Ƹ�1��5��
>X�ƥ�Z.�%!��U���#d�� @���n��x.�͜ı�p5����?<nk)�X_��m6W�t8�u$�ᄧ�N�ME���y��+��5�X�w����P(�~>�vZ�#�	|R319�u+����Su�1K�,[� ѷ��b��q?���V=���}h�osd���گ�TK���C��b���;���?��U :�����ˎ��.ѾfA���3�?���]_�m̠=�B�,��,�r�S�Er��t��&����8@�	 lM<vB�kΕ_�{^V��.�V��N�=�mW�l��B��B;��[{2�>$�!���IwI.B�_�5��	��ތ^(�R�BM�h�U���V��ۅO�m>���X3���y���+Ւ<zz��$-�=�)���bp�\��+Iu}ܦ�̞9f8;!�7�Z���n؋�?|�Ӛ�i�ӑn��>^�#�CT�2y����D\�Nt^F����]-�Er�D������x#,W��1�<,�Li?si�$<��}|���wkzAd���}R��.��ǉ�.z�L*L���^f�?>�0�	k�g|�0Mk/F[��U*i�'V����������3�߅��To�V��Y��Y%t0b��
,�O���} ��n������Q~(Hs�Fo=~��ۯW��R���c�Ԕ�f����8�Ի ��`��]�M�n�q��ED�)������*1�w~>-
�����Z�m�<k�<B��ݻ���Q}����᥋X�I)�����H=]��+.T��@��(���:W�/l�?[=!w8�6���]b����-LB���:N'��!����߼�j!�b1g���p�����y���'���i�ك�@uVQ�7vcP9�A��f�m$Z�f=����+X�l�Mr��_��c�r�XF���.-G�i���V;3�xL���j�=���Q�D��e�A�j�&�\��T��s��L��:��z�~�筬�bn�^�؂�.a�vݲ�`�Ƒ�����2����������'�O�ȍ'H����";��:�'�r`2eR�{����9{��א\����n(MWҺ�q'B���x�H����n�Y�+���M�;r��G2�ziܝ�����c ���
��a��y}r��ҝ>;]�h@��Gy�E�Ni��3��k��鴀~�P����㞟�k*��B�9������o�i�bLW�m6����}����͟Q1I�EEҸ��a`�`���b�͔�P71F[