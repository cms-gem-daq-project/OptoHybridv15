XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[ڎp(Q� �J�ʎ�!������.����y��j��ΰ�밓zɅ`�>�:�א��j���R�j�%j�I��u��}ZR�R�D)Yv���17g��W>D�D;������޼��rf7Tf4;绩n���a�4"s��H����N�&��Z*\�&g�X�e��^�����@$���j
��do�3�L��S~����������T�%�y����K�mh��3�`7�Yy�I�A䈦8=Hʤ�D�΅��a^I/))Uө�'�-avS�t��G�)�T�G:	�.�I\��H�~ޭI�J8Zqr�������IYy���~__,����^/���/�[K�9"춈�k���]�ދlܶ"�	���q����S�@��Z��/�B������i �2��hFVpY��S_�T�?������?8dD�8�\��,r��3�1t�vU� [���D0�����mT����9+"�@����/������9.�EU�L��g�j��,"DH����J�wY��!0���.0��;�F��L�*m��W��Y)]G�3�(!��N�B �0N*�N�lt�n7]�`�q����/˂�̃��C^Dۖ�%3F��������C�xm���'�'��LZK��Q���ሑ ccX����Gw-�n���C?d�;��wʘ��Ԉ�3_�g�n�9@J��W������
�4��&El��9K{�t�R;��g(���yv�O�'��s�4f��^ťc0XlxVHYEB     b05     370�'��-~�o���o}�҄>�mG`%�t<�s��!ڗ?��X���L/ɺ\�=�ā1��6]q|U�;D	gX�i��R��."��F?֎��	�� ���Oɨz�޳��&��z:�'"�&&�`�U��N�a/z�Of�f������uρ^V(<����4����5Y�(�[��$&�z�x�s ��I��/T����}�x̒�_.X�#��ӟ��<��h�i~,�4 �H���r>��z�$6<��-��VQRTw �w)�9�\�wo�F��Y����p���6�	�D�v��=v9�-e��Æ�3r�/@���JN$�b�=Y��"5��t��h"w�����'�m2+DKs|�*&�����)	$�d���ԕ7��Q�ClBU��o��x�jr��M)��T��/
4�6Gg�^`Q
�~mV��j����:����^�U�c(a~�C���1�*��Av��榦����3C�m	2��2�Q�|�]��U!iX�2N[6����O��B$446p 6�ݦ�	g��YUظ�&0�������o��-�<�NQRɊs�?��R�$��d|�|P�5��a+�^��#Tn�J*5�A5B��~�fõ�|}S����t/�=G�)լ^�]|X/ɰ!�eO��ς�P�Ul59��"V��T. [\a�b�:���R0�e���3_�V@(��5�X�l[դ.�$d��s;�$��	�W���أNC;�ۡ�*u[)���<�l�EG��S���":�k�6�;
c�N\��ґ�$z�H�~���z�miX;0-F?E��#�8^�|s��awu�)0T��7���H�V!��ښ7xs�]���@��ٗK����E3���S�y������g�yG;����