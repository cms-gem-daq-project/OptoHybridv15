XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b.�s��fa)�@;iE0!�6S7*VՒ�v�Uz��0+bgؙ5q⠪��^ǙdK����C0֭h��򿘱�4^���G8�4~��9$��_�?�ʈ֘&���5P �S��?�+K踏�t.1o�Q�3i�$S1���I$��<�#(�#�OzFcl�V*rU=��Y�Af?�EՉQÂ�z��^��JSŞ�:cU,���� A,hlf�7�ޒ�i����!�fK�*�I���O@X�o0�V$�&1��J��%X|-C�]#�^-��Ne:�!Qh����9��%��1���B����TtmB�5�o�JaA�����;�!T���M�v��X�7�^I�Y�p�ґ�(���i�<�W���i �I/��JN�����t�P@�x�0wKG���v��x�����$id碬 D�C�Q�V�H�B3m;.Zߘ%�I됣"J��H�AA
����9��w�� �.����s���L�⿽)��&JF��:��7��w����7���W(1�k�N��4�����{�n�b���[��B��ǧ�i�;�� ���O�ƣ���~�H	���ġ*��J�u%�#�l["]�A�K/��M�/o��q<��cs)L�[-���r�o�u��*���7���::��bWk⣱���7����4�d㷥�2���$��g�����n�*d�.��qH�n���q�sն�b� 1g%�u<z@�"��qG��j�$�H�P6-�f�I�?�^Qb�.:�cAM��XlxVHYEB     4fe     240���<�,�u��a��J�#�� P�,����ٛ����p��;��D�v�������=��g��^Z7�7���[cmL��}�Xm}&�v*9BY�hX������<�PB�ts�Gb�����G=W`��2b�W{i/�I���3�l���tܨ+�U	]뾋�FQ����)�)���� �=r`Ԅ���q��΅ě���,0!�;���e���LI�RQq�����Z~n3���،�u;b��ֽ�F�kqꌭ�'/�/��`����R1\g��7�2zV�e������6���L���t�-y��]�
6_:���қb:��G��A�����M� /Z���0B(�Dd�A���|f_�?k�(^ �����ֵ�KAJ� \z��h�W
!3� ���v�rQ��!�:e��7��)8���%�Ϟ1b�_�B�Z�Ux���ۑ&6@���g O(�ꪬA3������E�#���tmvs�֠�՚�Wd�M'�.���а�U���|@�7��|�l��A���^�����"���Sj�Z	�쮠�l�?�qr��k�X�?t�V���B�