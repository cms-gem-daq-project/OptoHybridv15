XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�N�o8*j�Btj���v��VF�S�r*isf�&N���Ym"�qx4bǩ��@4KH��@ոޑ�d��T�oѨ'��8�1*q�u��\�QT\7_��zϩ_��)˛4��*��n˚憕�����>va�98fЄ�
�bO��ʖ��^�Gr�6n�ү��mX�r�.%Q��Cf2���/D�s��Cج+���l�������f	h"S,�#;���X���$�{�e��4���@CZВ�����<��l�5�a.�z�(y�R�$������d��Q�A��d~>����q������Y�1�|���T��#tԤa4������\/͉:��>fZ�\�az��%�)s/�¢�ݑ6�I}��~�T
I~[-�����,)U�)����0B�J�К����2�&Bo}f�ǻ���}֊y���p�:ǥ�g�F����Yk��Q�y��'	?
��r_@rf�]�-ַT�z�|�Z�vd���gl�(4{Uc1%	D~{-��mmU1��<v[��_��^#�q%D� Z&i#v�.�e�R���]��xe����Pxf��E�H:^Th O�Xە{�|h\�-�v�3c�V+Pa��~��`<-�ȅ^���9ыu�8����$i�1�$`vB������د^��x`nj�0LI��?P�{�WΗ[��6t.�8�����r}w�+mA?Wq��O~�;@|͏�k$���Ԅ+�酽�C3*~M
��5P�/ ����\��t�XlxVHYEB    8625     ee0t2��2<  �YQ��\^���*�&�w��e=����~�T�^���%PGK$
��
�ۍ&Dzj�} �Ձ��.x+Xj�S����8	�ᶆ���T�o�����Ju\g�i"�Ŏ�������?�FlHd �+�ٓ�2�,@����BpVp,9Ҵk���I��7s�ښd��a (Z��"����(gN�h��yb/�O-�rs����-Ts�p�r����9�j/��s�ދ<�Ѭ#�u�|�ꦈ��6i����2�j����®A�Ou�����Ms����Sa�ƴ�k�3�/ �)ƾ�&��5k�Iz�V�o�^� ���=���������~ϯ��tI��y�G�X���s��j�ҷs���O eYrc/Lf���hl��;_��>��a��=�ѣ�)�7�ր/�sX�~Ȃ�#����]��a�)�w�k7l;޽&4�U�T�� �Ӕ$��-���`��I����H��},�4� ?}A3ԭ��O����=y�
�[/���Dj�f�{t�80�pY��8e#�f��o����R�7���s<pe���Wl_�����
������ ?@��a�+\�i�����w���2�XC� ��(9q9��6�Lxw@�9�I��ok�Z/4E^`4Pެ��Ocʌ�j��wV�>�[�^3b4:�<�o#P͍A�V�Ԛ���}��Ʊ�z�'^亨��SM1P�gJ^D�X4�!�Eq�pA2�EF���
�\�wvU�v��wm׽�'�1($���Y����>'.��Z���%x( ^B0FUs�b��*$��9�[��0�N��C&��'6�׮=�����K���x�@�q���<��l@j����gͼ����0W�_e�����ٞO�zx��T�e2o
�bW������6�ǖ��� �������zb(�_���csa�֎�2���c�ì���V�%���F�Z����@��*]e�܁&����,�Cb���C�9*sy>��MP(��<���s�uQ��#2w�f�����r���$X�5嫔.�"'��a�eI�ə�!1?{3�9	��4����#��չ3ʨ!��y3aM��:)�z�qԒ�T����d�뿅�ؗ��x�3qE��i��ū/,�	�|t����ŧDc�FHDs?�����{�k�#�X�E13 �5���_�ߖ^G��Py�BO�(��M~�xȄ73����$_Z�oKǘ����א	3Lb�})$~H�ߖ�=�t-�i�E��s���󖢖6HۡPyk�~,!.��W'Y�F����\mi�O�3/!rH�f�?�J����7�ָ�$ w;?��OJ:/�	�5�E�*���r�����5��2�Y�NO��%�B$t����7�h]o��K�E�O�p��0�m]�"j'f\]x���:�{�1���J�����+�1�hZeg���W�T˼9���߹P��v����г�9�N(���!4/�=���.���YQ�%3�5����櫘�&�@ݓ���T�@��vX�fp���@)��q��g6<��Zzt�酭=��t�TC����0`Y��2���R���tc,����
Y�!�`�3˚���[����ו��P���e���c�NY��Wڹ�������D�d3%+�XR,e�@�?Xzr�\��w��n<�dJ�݆�n1O��$�O6e���o�����;δ�k���8�K��:	�Ho*af{&��KUȃ6�2
g�vr�^<���1�Jpv�86v +��ZX���G��l�b��do&��Z�K*É��ɪ�sn��Km�_��;SW������وڛ7hR1
�cU?��\�]�N��Cw�q�%�����A3-����?a��_)*�i�+ ���Y��\3b�7�U�S�Lo�u2Mt����6���T��Vf��oa��j�f��EBe"��Ȏb�9����(�&Z�ɱ��=Ո=��Mmk�z������S6-�4�<>�$�.�y����昒"y҉ȱk&i�����ߵ5�I�#K����&�4�5j�E���RWr-N�p�{�^:)�����j0�%�䘘M��|���"L�ñ	�*�_<ܑ�B�Ş"͏9�s�$�a�3s�Iڿ�N�/����o�2�o 
A�h^)1j���5���4��uS�W��(RM;����G%T ?��Eh��5_y�b���/G,�EKh���=��3����B�U�p��q\�K1��)K����W�a\���ֳ���E^�Sm"̋�V{	m�z U-��#�W!�b���=��;M����c0��AZ���:�-��s��r��m���2lͬc�sR��>��i����>vm���*p	io��dש��p~֞R�JzQ8��Ǥ��v��9{�*T�*�:Z2�pf;YX�i���w�V����Q~�э|�;���$S ���`�����1YYg%"�l�U�L�ާ�@l���1(3��z@��v��2-���Y�C�}\�9����w���?�o�eV�V�
��Xa$b5z��?Pt�֍_� )��m�J����ʪ$���%-�dL���E5{�J'V�6H=��i���v������r��17�TT�l����<SZ���b+�O�|�k_ ���1� 
9�~n�~B�iD�C<��t�K���r��UZ݀
�(���.,dp��>X��D2Y����"	d�L�$.i�}����d��8�q��-	��L�7a�TĘ�O=%؜��I��8����"j5�u�q��8RPczr'^ou؀;!���<���A�y�2!}���_)bBI�V���z	�=ܜ3�`a9�I����ɯ~��g�hTq��2(��+�X{�����Q�U��hL�gj��_��;��!��XX<C$�2H��I�h?�i�L�h5M> 5 ?]�
�z��@R�2�:�ٽ�m�n:t���ą:S�'��`6�&-Ÿ��D82�L���{	�5M�PR�a?d����{��᣼�� >�k:�m�a�,ʊM���^�-h�(�<6̍��в�d4�a���Z���n�˃FV@��hPX^�-��ߣ	�4̶��b������S�)6r�Oi��2��I��x��>�/u	���U�jT����#�Ι��mA�a����Y�w��L؟��J��Z�ea�47
��S����HA�I�j��@g�F��t�0�ِ�.��hkT���N�`o�r�1]14��kx`{�<���1���y&	"����`�(V�!�^y�ű�IUn�oN�Ќ�I�
0�!��hV��<��8����u��(�-q�oe+>��CG�h�n|_V�8R�Sn:.���IV��<)(Z�T���&�-Ҧ�5�$����pj�)r��^�pa�iN�5�[atdm6�^�r� 4|�@��G�H��Q���)�� Μ3D-���[��h|1��|ZSl����O�?�Xb�g�Ll�X�1����V�Oj�U�8�ZG����z������-..�n0��S���w+�w�P�YDE&Ėh�#s�W|XӍ�z�c�
���!B�KS��� >��`֓�U�)B�Ƥ.�gL�^�<Ux��:��$�FQa���1xh���R=���WY88�r��D�P����0=�(f���ǰ��x�c�����H�O�)<;��=��o����p�ejz���g���FkqZ��"ō������!NYJ�lU������yޔRf�+5���3�|�pB�.�үk�r��򺿺U�j}M;(���v�