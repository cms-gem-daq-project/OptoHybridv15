XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x��^�Bt�g
P{䰉Qr��ˠ������/��p;Z�����짴%ph�{Ґ��<�H��+���B+�����ΗE�h��wi�������;��j�DM�6�0��S�������r��q�Jv� �?�3�ͅ�Q��<�/�� �4�xv�M|j��KM�j�F�1��}Hް��L�=�ԗ���ٟ���R�y7�vn<֑{x~Ϛ����$<�md���ݨ��]H����u[8O�{�y0n���|�)����}w#���Rp�GK[2��@@һ�������A�lgO����uih}�|u���5��5`C~g:�����B�U��J,����Ҧ�&�����%4&ru���1s�_}�	���'Q�E!�ÀSTc@��%�Sk��B�,����|W�xhU�1k�F�m���o��W����_r�s�p A�\��a�8��/��+@e̝G=Z��Hh��_	��D-G��/G�n]�]a�/<�t�dP�a�3.��UR�A-�R��!{��������~>�c}Dtk|��i昃 Q���86��Ͼ~�.��Ο�ǘbF��Ӿ�-éU4ĈF�]J�8a����1��xs8���c�KI�J��d��Y�Z23�M�hg# \��J~�DW���j(������SSκ��:� ��)����f��Լ������3��G�u59u�~~l�:⦛vh�S�,�j�{94B&"s�;�����HZ��D�j��~�W�?�`p�X��/XlxVHYEB     b7b     470�0r!b�Km��ɝ<#a��m�Z��s	���Z%̢<�6�?t���2�q���i��}�����8M0y�I���"ԥ��Lq�`�{�:�}����v�ͬ%'�ƥ�kbb��rٍ��|�"x��7;�0����+����G;Ҳ
2ɲ�<�b�d��<��d�����5������%��2�˓�W=Q�^��m���J�7n�9���ri �� P0���wlT_���G����=�`�$�Jm�F�8)���i�vVfj��$��C���
PSm�3pylq�E�u�H��@"����YQ����T@ ��8:#f��0(�7�+����M/�oi���䷚�1o=���^�<��"�b7�
��z��v+�ô�]CN���ҦW�ǭ����^���L�MU��'��u�`��6�0^aJ�����u.sN�j%���Wso#)��(����Xع�Q<Ğ@�n���.��L��[w�)Ij�J-�1�w�����Z6�c}���h Q�$�UF'|�u�01s�A�eG���չ`0����Htp za�	���1Dҡ٦�fL�4B*O� *���rX��T�E��������~�5*@x&�6��iSD2��c4~ջ:���mw��.�P��:�,���F�7�RKh/�tN$ �[KZUV�۹?;�I���T��5qp��X����ȹX0��ƍ7�|u-��t>��'@:6��x�XZ���6ӳGi��a4�--D �F�=�����'I��>����Ն�uC�Ԍ���djQ�ƢR�E=�q����Ry����_1U(Pz����M��*a"�Y<݁�7��̪yU" -�A��qQcY�r����l'YO�ܽ01������R���3���veҐHѽ�3t�Ƀ ���K��cR{E����T�zQ`ӑ�n��t�Gp��Kx��H����C�ya��)�A
a�
����i�Q�A��%#�~rJ��C�w�M���/$c�:)t�OU�Z��`���Ie�F���PGr~�0��	#�~u/�;c����t����A�,��fҬG���_����]p�2D��.���S%�����T*� TAI�A�˞�q1Ibg���