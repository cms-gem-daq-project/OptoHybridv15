XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��} ��R
.SW�(A3'�v=����t�ʋ�w���ό?Kgd҄NB��vVߣ@��m�8}���ׂ/X|��?z�8�]Ja"%�vCà��Y�a�:M��
�<�nM/�>�|�9��)��uϑ���,΄�XTd�_�I��h!	��"�7��u��Wci5��3������F�����-fHĶC_"i��+��o�j"�B�gJقIފ@�b[�K�G�bv�R�2���,�Z��������7k\R���7eu;_��l)��X����X�30�Xp�ɹ��/�i�� Ӱ�sBcu�@��*#J�U1RO��nB<����U�T���|�gL��y��g�9��������HH�Y�u�^h�>Z�t��ybR�N;u.\�Z��_���T������=+�<_���.*��/�!���)��c���a�D�{}�w�e�*�$sލ���`f�������x6�E���Գ��������<�A`��M�0Z@�;���J�Pl00�5WRO�[�A��Y����^2��(��X��O�<|�ؗŉ�&�핸�� '.����r�RB��H�!?ߘ��(E{����Vm�q��,/��	"j�1�~�����n0�b����`�
Ԉ����yܝ��̝!0�ﻒ����=aG$l�YM������7��rg�	�������:��D�E�ʞ����?��F��}W�>��+1�����!g�p��e��c��Hz�HFXlxVHYEB    5ff1    1040&�Ǜ�C5Qc���/�MQ� ���3D���N���5����(U�l
?���.O "�Twt��RaR�U�{�ZH�CF��c��2��� $�*#d�dhD=>����(kκY
5��/�"
͡j�?«��@)yY��`���%G-�y�c1�H�O��C�!#?�r�ɀ�R��hL�$ƒ)��a D�ߕ�������8����
�,f�eS���1��o�h�_�IuQ�D�_��77թ���Q��U�κ���n��0׀�D����Y��ه|k�&)M\�N�~d�C�%���q�3l��x�����vj����W����:C����W���'�9$8� ��'I���8_٠z�[����XIt
�m�h�zfp�m&cٽ1�SŠ>#���P���n%�Jܺ�wҜ�QA<��v`��+���^z6�P9$AH�9�Q1����\J&����Q���I�����U�w�I�+]!:�w��a&!�W������Ȕ�T�b<��L��ba7Os��x�y�����E��-d]h6��D`	R�Z�7U�B�S1%^$Y�I�2�I�> %BĀ�|0x^]-�#!
,mk\?�XN`"Z���^�[ ֢�R��iYz;�T����k����i�͏�靀y�y��|�� ���U���ǝ|�&��t\q�"�+��������,�W Fb>��FJ���Cg���؈p�-�g���I*��@=�J�CJ9�=g��7SS��@�?ͨ�lS�:�wxJr���C����l)�qX?���<�4f���g=���B?Q���Rg�SXc�h�"��#��O^����r#QI.V�T{�;�����b+D�4o��8�h���z�)�WYMZ��-BKߐ*�Rs&�(H�����w^9<�}c�� ��I��g�"�]1ipth u���7	�>x��[��ïjbnՖ�v��S��C�̡�8.����K�kp<N��.�q5�W�Av��΃[��}���a��+�Ì�\��d� }֟����j͢SAڣ���GD�Tj��������W�ɑ�"r�����w)�h�*n�.���b��8���yV}
m�Ҍ�+Ls�Lo����C@`�5���Ld�.��.�C1⅟��p�"\,�ԂZut�v��?��U����yb)�W�q@�j���8"�¸_<����N	V�G_:p;+�mO��6F�{<�׶Yi��G�16&����� �Zo1�EgAZ�55f]�]g�!�X�=#��2�0h��Yg��4o%��A�Ӄ�@����3��Z��6K:�;CI��3���x̓��yO�F�,j�9��V��ȥ�s����!$���6�[.�褌��<[��/����"RTJhu2<X�$������%��{�O�+�u���e�Ȯ�r��K���� �(B��uY�m�;]��z�yBP���:4�	�M�<�q]Qm��QDZǢ�.�i}ݢ5�[��:�K�M�����$)32�~g+�u�ŪM+fOaF�B���Ӯ��C�c��<��@"=sT��x2`	U�Af�
���܅<� ����[���bT᱄=�z��]�`w�ȕ�1j��Ղ�:�,mK�{N��6�Y��S@}!}��X�JD��LpLg�c�|�a$�]g��m?�|Mb��b�	"����|O�����[�J��b,'�gy�}Y�Ju{*u���ͻ�oo`�jUp76M��9��ʀ�:F���X#!��`m�,�6A�z�c�W�7�{���jp����MW�%K�"sl<�z���a�Y�_�i�A�Ɔ�V{��5�B���l�ֻ�Be� ,I&l?�%��k1EXy�W��8Ԭ\�'�GZ�t�H�4��Vo�<f��sHo��A%L���mL���A�����̀�?�
4KJ��(r����*��k����P&x/]u�g�M�hN60H���9����_y�l�T�� T�B����N�GKT�}��X��o��ѻ p�S�~tI�~���tҁ�10����3��ry��CBؗR�r�����:j3�����E�{G�~*��#I�ahb�G'��M������0E*���O��lw�r��䷸�<SX���ι*�@�R��H�Ý�t�����0��6��C������J2��.JV���jRL+��Jd��L=���\Y�u|�P�#��oB�}V%y?j�4�Mƿ�Dq��a4(��`X>�
�ë��z�T�I6H�M#���h)NY�����5����#o=��h�����P��������x'�m9��@>a{�;�$��_�VO	eW��9�M��m�׵u�H�h�X�Q�J�Q��+����~�\�q? ��N]��U��X�J� ۖ��1N�k8��BC�uG�7��Z��0�hp5����X����j� x'�(��*m��������i½"hpm���Ěw�֜���Ժ�(�i�lD@��~A��b�?a�g����2b�Z\,ԓ��5�ȥ� k!=B��̬=���k�*=t6#��w��d�����2���x�PÑc����.�U�:&�h>l��0��I��˂XT�IA[=����a������|�l��<M�_�q�����2�:anڝt=^k�
7�T������y!�'#{�۠�E��9ȁ�mMu�������\�]b���M��L��x(J�L��#�o��u�,���)�W2���MAUS��{�_j�Am���U�䜯9�;�L��TC�����Vl5:Ϩ6{d�sA��]>l�i��y$)�Wm�sNI	Ow��K�&,�jf�''LK_9�UN�&�#Ϛ�oM��ѻ�Y��x��p
���U怇Ŗ�	�7i�^
{�$�S$yŬ����9S��ҵiѹ�̗f��!긺'D)�G���
�4��O�\U�jo���h� o�5ʥ�Ǌ�%;&���g%����ke��Y���x��� �ȿ��������R�ם�G�/��9*p�%pv��T��~1K��i;�5=-�wrjo���ށ�����Fdh��������pﰛM��l�����5s|)Sa�I-b��Ǝ�L�l�R�ܨ�~gWwU���5?#YBPB�߫���'Տ�XZ�t������u>�q]�{̻Ӧ#G3��R�2�ϔ���K�T��A�!��ո�ܟ.2�7��
|��\J�<d�w�nA<%*w��;���M ]�"�/�4OU9Q/Ry��\�\	�SLy3�*�Z{��Z�y���H$'	ُ��2A�MFjbvpF�$Q�נLP�W:a'�Z��6��u��֦�o�Y۲����
Ȁ�
\��X'@@����ȓ��J��6�RcD���K+n-�<u��:���x7n���,q��d�ݣ=���7������fS����%9Bx�8�bc��b���y���T�-���g?*� S��m��� ��c��Z&)�P �y9r� q�DDF�tww	䚨� ����؟��P���m�����R�՝�؏3^�`! *ד�k�6��œ�,��u�@`|={��nڽl�+"
�{�ԕS2���-��<&������
���*t>�5����W�����Ŕ7�L5�\��Hw�.Lp�
��*;�g�.�Ιuű)4�8cT/�P{���D_[c�.l�Μ��JQ��ͤ����/Ǿ[�k%�d��&�H��X���t)���	�7����>�^�EwBfX�q}��29	i���&�[t;�G���6Oٮ�������H.�h��p/�ῶ��w�H�������$Ym?����,�l������f��"���,B.Dِ�����;��@���g;{�V�Ѱ��C�es��
/�S:A�r��2��\�xE&S jLCV�ڴ��#�w��|iZg�\��.��f�g#lЄR��^��ʍ3>a�r�!	�>�i�D�&���V���q���r�}i�5�,P�T:[��dJ��^a�|I����1B[����s�b�n&,q�N��&c3h핤�ut9�p7��N����U`e|k?���qt�(�ṭ^�g)��s���E�w!?� ,�6b@��l�� �'�-����ک���