XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W��b��ceS�ٴ�<*��O��($@���Q�N�����P'A���lC^4�c����R<���Ws9���S����Jg����]��ccSNl�U�zַu7�$`@!V ��-�Ys/�-K����d���G�W_Ǭ9 ��,#�I�Ә�&���
�����y��lag�GNb�x��q�8�NS��R��uGI�2�2�.��R�v�y?��6�����SY����XD����K`5�tx�a�9-Y ~,s(�i"i��'P�Rꯣ��Q5ə�B3=WӁ��2�f��eR��_����g�@k����wY�;)k�`���m��X���j����������������Z*K���	0�w��ZL���ܳ�y�i`�^�#�x�����34c�4D����V̞��*�A}��9���~K=p�I�8�#��(3<�jЈ�(���:�M������7ڦ����'��+�>�O��"U�v�~j?����/�j�Ը�u�>I)`��Ǆ6�E�p:��!����פG�vi��;��YW�D�>v�żAC#.ߘ�p���J�q�y�̥�X�V�����ɌM��U_8X9mD�w��RZ"wο�q[=P�y��<��lI.�9t`�u���|�eᐉdsӢ�BB��_V�|	������*���mm7����	�7�Scv�>��F7c`4Xk��	�e���Prr+��gN���Jr0��z�;gȨ���Ue���újn�s�VT������WX�~o��Q7���b%6@IfXlxVHYEB    1cf7     7909]}��O��"Q66q�)���#H���"���D�6����3[ ���г��᥊c�Wxr���Y�g�3
���:�s� �:��{�/��E�]�4��K�����ZM(@bē�)�9�p��˗�Ӥ�W�O���T�?DG�X������Ҙ�qN��m�E�<��55�6���Z��Z:�K-��K��3�������[��g Ã��On0�D hT�z��HM�fXH�#��c;Qq�>�VͻV\��ck	���S�9���S����!@zch��"����Zګ��#���Rϝ<��!��z=�Mo��T��?&wb���]��+�ו���y��ƌ��IBl|~W7؍;5V���E�9�n�X.I<���3�-��n{�Tt�><D[���W6$�6�h̬$wNWZH2l��48�n��Sn�r��8=";�
�s��B?=;�T��د۱j�0I>��u���R@�%���18��<B�|X�� �X�(����ǂm�W��B{((:�	nn��b�B��%L�i���~W��0IF��^��Xc��!1�J�iV�ԍP!jU4���]ՋKn4�Oભ�s�h��/!�M���<�
'���޶�q6]��;�T/K���>�_[S��d1�z�'���PQ��N-v��0�9H�X9����~���w��=I�$0��h�V�O2-��sU� �+��q�K+\zV�?|�zɰ0���1��A�`FJ��&Bh���6!T)��i��)��a��ʛ��ȫ��u(�Z��5�h��A���u��C:l�b������
�+c��A4AQNF �o�=0|��=ۿ��,Voq�>�*iP����,_��j:Y�0&gR�>���x@6�S��Sst��o�o�KB��z�a1�iD7X(������W�(W�_x��[�`�I��rׁ�4����S4T��U���}l��Dp��Ag�Cź���d-$��L������&���1i�fW�Ӻ=������Fm����^�y����y�1���
}��e�T�<�3?���r.cш��O�X�ьK�{Z6��d�H��$A����q��΁Xw��Yw��A�J�5h`����)�������.�C�r�v/���`��k�^��k��Z�K�+�#���lnx�-�*�T5�k����K?~w�N�Gj|���5����Ry�0 �s=ⶅ���3���w�S�?Ŕ�M��� #w�\��^ʣ3��I��C]qnPb�#󋻛/���給/������"%\��r�4�JW� 28!�[]hT���k�P����@���B�Ȇl���\߉rs����fŲ�=+�R�<6�t���A�{ݞ�l�S�S�)�H:	�b��Is}�t��J*b�i�h~�;��
s���Ă��m�����IQ���PV����n�M�$������3ٔ�$��$����s��N�"�^����i���(pJ�o����d�Hݐ��D�����/�hty���ꗚ��ʹ����S���(ˈ��3�@7-=O�� Wt�(�X��/�zR2T��WOoX/}�\�I���)M ��$�j2�I7��7�ryM9� �����Y�NH~��L�-��u��&_�/�h��g�@Hc egf�#㕇 �G�Њ$��S�S�s�m���ö����o������P=CC���L��^	�X�3�L��"3�yDZ��Ғ-v������3��:Vb�:����S���9��>�Y����KV���}���%E��C���6�xIM��-�������Inr���.b����B3=��1�vZCԢ�v�;o���Mg�n��;��4�tk�E�A�,Q��b?TK�u�3��OB �q�[�׀��e'�&�;y�[�'��S��