XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`Z7����@�''b�� 4֊k ��Xz�d�<���px� �e��� �}t&�A�.����_�5���M�)�PĻ�Z���U��׃�nR�(�)
>6�JЏ���j�/o��:#H�DX{�V��uZ���dX�f ;�&C�Qg��$�eZ3���ڛ9���2���t�l0����
����m��Z�1�w�d
�������ޕ��!�r�ƺ��(WV�i����r�4_t�x9���G`��yx��Ч��.%���ݚt*�Nn�O��65�����ô�	a�Qn+H���!V�(��	0�!+���e�7���%�PY���m"u��Y�.��'�����MH`T���ʒ�kW����U����{=����0�s����C�p܌�*B���R�%#$I��w�Ǉ�K�h:Z�ٛ����!/ٍ�ZUJ�6��K�<��kǇ�J1���Q���1�c�5xp��ʲa�Y_�ӈ�_>�H����WJ�s2�W�%{?�mG]\�M������w[C�U��W�SܬDܣv��Y��@>.'�BN�L���f����?��	�/-!�;W's^�X�}�\v���r:���T�T��h�I�I��ev�qF]�w��O�K�֒7%F�h���I6YJ�ai�$�?`]�U���6j�)�)(].�x
M���fL��2Q�L5�2>u�����ÕҝAV3j������!�7\��T�p�iD/�߁II���wNz�͸�XlxVHYEB     b35     3d0�^+��63g���<1�����ro�qj�<l��`�b1����D.V�c
(&[I.�&m��ᥟ\q�pwL��GT�f��{	R^vz�+@� \�d�~�n$l�	��a߻�] �Z��i���z�:��ʗ�9�~�ɶ�͋;A���G��s�;`gߐUЛW``g~���w�{��N�&p�����浴������L\�jv��ge�d���A�����_*��Ą��$�I�U��kL���òY	Ei�+��a�ژD*U�Ս�n�Z�)�"p2pM���E��v�V�^�B�t�"]�f���z�lfF�H�Xg3��]k�|�@ɱ���n�o�^�;[#�A%�SR�WYmiJ�{��{�\?���P���[�ʨ�9e��R�p�����S	���?a~���q���KW���7D���p�&wg���߰��3b\2��n2TK�c��c�����h�Lrx
�}�n'TW�`|�eD�I,ZVSC>b��ewb@в����;��#��![LCY7����D7 + ���N��8����LeF"2
]S�^:5��R���m-���hA6�XPNr�����<���0?!>n[�&YE����HJI倝��k�5Ϳ��>��%F��mi�Z�S�����9I��ڨ��E6��{Ot�J�Q�+���i��o��F�eEU�)�.�}8D�}����լnٓ����t��p���'"��a� ���BJ=h9���a�	�m�/J���9�cŬ�ӛ�� ʌ鴃��|J�..�R��%�61Z9Q��F�&9/d� Y���Rs37}�mdT� ס�F��&<����D�9s��;��G�+��efxq�W��18��2��s=y���_MϤc'?�����2�{-����e�^8ӳ� �a�:�faI ��\�r�\��ʩ���mZ���'U�\��Ĥ���wح�)�P��E