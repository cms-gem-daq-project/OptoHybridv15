XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&t�������̾��F��,��@L]bw*qs��:  �� ~jT)�,�9�����b�����?��`���$5sct�N� x�K5b�����E���;M5�M�+�i���Yւ������/(�%W��yQ_|R9ѧ�+������W�g�,�mQ$m�L���;�3�B���<���X���zl)��TKN꬇�J��-��!� :sKu�'PA6զ����#BBA�W�촁q[��S��8ґ�R����RQ����S7�(�	��d��+DFiqd<��n���q@pb��b����+\+t��iLi�5���*��a��`r��/r�ڏ1��!zXՊ$�#��pa�3���a#]d�|=�l��Ll��y�&��K��a�9�"}��Hgɑ��ԏH
i�}H�ǟ���W9������y��m��/��Π |�S.��i����e'���l�4�o�`ĉ�� ɓ��x��P�f?��Kk�s��5���7e>����H�����6�L�ɻCj���k�����o��d�'��W���[B�f��b�~kD�B#�,������d�7�Q��0o�_U)��IH�3RG��t$*�+�QNʄ�P�00��9��(����%�Y�!A�1�r��ǭ�.*\��8�~1�CGIOpc7\�e���+�*����P�ť&��\��i��K��苏�Lgo�?���\��V�%D�b�+����f�&���`�k[87�u��ci�'XlxVHYEB    152d     5808��o�1n}`�?�a���̵T�	��F�'P��b1�2��@`?�0#��%f�����b�ry�&��N���d^����Nk.�N�"���ʬ3~�q�IG��!+�Tk���!�,E}K �ɠk禣=�;k���[P`A�
�;������"��F^'H��^K[g�H��j�ۦn+j��m�c���*��D�8R��I%
垣�7�#���A�(�e�y��E��d"��t����ہ ��D�����K�!�ҭ �� L�A�$8ЮR�#�߷
�U���h�������ti�3Y|�J,D�,Ջ:�"��e�i����2Anu,�o�dٮV�����Al���g���E�	N��K��?Kn�=P�,`�:����#��8�`G��樨^��� � X��r��0��e ��1۵b���XR�-��%�hӂo���e�M�E��V�c�]`��P M�9�,N�T���?���#�/A��x���"d{�U�?��c�-h���:�B��D�7�AR�7���R�D���k5"}�����F�-p�gh,"_���Kb��E����.#ō|8��TR�
��{����� }V)�œw'�p��,�����c�!�!*`�S�T��#���oT��2 !p����Q%F2��w�i�� �1�`)�`Ja!����ٷ���p�Z}1a�7��f�	H+��;�x˃��(y�t�t�(S�}E}|��Dkܑɬ�6r�=���L�v+�)2{�CBt;�#����������cɹ�Q�48m)�:Yܨ�AsT12!/�i��Ƿd�y�����2�wCr���y��z�2o�/���Fr����|K� h�Ai�0�����Zlgs���u�BY�F�ä�k3�G1̴bTq�vPCo'Ȯ��� ��j���i�׼ͮ���r�;l���R���锂er��jpm�g�!�fP��rVuu�j��^+:� 6O
�S3t
�n�T�_.a��Ρ�_$�}
mm�QJ�ΐ��E˴��w��}n6a8��Пk��SA*�C9����m�+ jk�r�����bn݈���	�xR��!���,��OVAB
Q�y$I��-ͼ�2m	���V�G�s>����Df��"^��$٨��r�/d@Nj� #��껝R���k��l��r���������ַ�ܢq+N�y���M��b|W�����*J�b�D�45�NN燋��u�e���,���fMx/Z��,l�uꖻF rR@[��
W�䄈i�n�|Ϟ]bR���!
h/�����V�^[ʭ dy/�Ѯ�=M�3�\�vM�f�({��]b J���˱oa���z��!��TOx��EG�çW�a�%��,ū�\a$�1�!H�긙_����VKd8��k��yA��