XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	ncs����i���߹�T���e�&���ank��:҉R�w%�,x�u����t�Id>����N����N[��K |qL�Y]C����K핏זVm��V^a$���?d3�1��!�u�"�#Y|�m���s�$�k?�f>����<�r����=@���=`��U�L� E�-q%W�2L��Q��"��m[ǡ�s�W;s7���Qؔ]\q��w�'n�:��Ɂ�L�L���&~Pɳ�%U�&Ի{�V�,"<~���lmN5E̹��	R?�����ʅO�B����U�[�G�E�+A�y���ׅ|�Y=�
,��|\JbL��x�>�KbkӶ9��ȳ؇��U�HSk�]���h�@Ql&r����M�`'!T�b
��T����j���j}�R�G	 c|.�@ ����|�\���������7�����Qx蟫�2O~�u ����P78=�O=��|go�݉�cX�l����$�C,�,�X}�߷g2�����i*x�S���sN�6 j�u��|�6x�34�&�.�_r�J��{W.��x����\�5�=ߒ���3H�Z�X��і��I���^��F��/��ϙ:�sIP#�c�0�Ey�z$v'��#���x;d�����N�OP(����@;�ಽ!9BqO�k�%�Z�1��H*���{��H�1���g�<�hp��MsS|�	^�|qA&����M����B��C��\�*������+ҝ�yDi ��t��7E߾�g��XlxVHYEB    5a4a     590�Q)�1�_�"��&<���ޠe4�~�����N�����RK� l>��@ׇU��� e����\l���g�Y ɾv�{�#%wL���_ I� ��0��u�\�Ш���Ϳ�p���:���OU���jW�$��mR{6��l�RvVnu�m�l�Ĵ�B~�@�.{N̻���p�>��I � E]�0=�B[����,���>�`ٿ�y��A7$��m������
s�˥�(�>�G���E[�>>o�3F�C�.��@��̣���c��9r`�pϏo�D��� �����~#�h3+��%�2&y��Z�u�nY9�7!��$n�jp�DC3��));��[�2tW�s���sL�Ƽn� �i� �i==�9�sM{�.*���S�S=�qw
@P�P�"�}Wv��������x�2|f��]�Jo=�%�e��,��p�;���T�7#�%뱵�Ҟy�"��[w��G7�u��MJ��,�m�}���9ztz-?�T9�a���Sre��Q�3�.����p�0V�4V��M��$��Mץʗ�P_��������r]�G
�Z^�Ⱥ(uB��b�f�P14m�K�w����Q?��8δ�$^��*�Di5;���sB�ڞ��3���ʭ��?u#R��:�&����l6pqq(��%#�P�.��,kI��/�z@"䯭�$.�)�K��� c��J���|��0G�ኝ��S�f��,r�
=�&7M�mc�jCPq/m�(��oa�Ĕ��]�2w+:S�<W�z �?r������y��_�3*��qP�K��{��Q��X� ��]+f�Bһ�e��[j���TU�x��8޿3���ۈ�6ˈ���^-��)�'G�<�T;-Wǌ�k���r>#�<0���� �Pʍ,[@=^����Ŕ/ֽK4��#�(���̈��}=�8�[q�-�����s]�殀����b��q F����ҥčh����J���#}@6(��+e�}�b�$8�a �ˑ�~й]l�� :ް_?�))�{��PCƟ���.���:9��e�ɣ�%���)�z��e��#�I�D_�h�S�(C����m�7U�0.��	�R����f~�L��Nwqmm%�!,QaM��z���9��ʻZ��YyK�����{ݾ#.y0�N	M�Y+��	x)���^��.�q�s���q�����a+QD��'^u���������3g�@I����)23��E4	ޛm�:�Cg��}G�t�-2G�˃x�該�8!��y���6�%���}.��r�mY����k`��Q�8bN���NC��>�I#��8�uϮ]��t����t�+i��'�t�j�.$DA�潠ʄ���";���}�)��0��kڥ_{]|�3�h�����<�:�e�"]EL�{�0�`\�X