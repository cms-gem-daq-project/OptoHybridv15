XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/%j5Y�l���Q�C�轛'1R�`$���x:iM�U Ek$��9PTI��V��A���6�C[�Z#�NɆ%�-T0��\�6�A���p��;���z���9����Sģ�3��0�q`�=VYas���#y	qo�x%�f7�)�^�Ռ^w{��<(�)BJ�M��m���'��&���]!5'ʢ����&C�eG�b�9�����E,R��_D�Ǔӄ�d
_<r�Z�1��ޔ�ul��V��2�LlV�-&$�^t�1(���g1�r��F:e���}ND����Hk.*�rq��PwVʜ��s�߮�C"碗ft�������޽��v�z�./�),SA{?⢷|GkԬ�!O,w�U~��L~
V�RN��w�m����?Y��Pa�眞�9�+.�wl �md�{�Yur�P��1��o����E@
�f���½�)�R��E�R_�.=FZ4��M�a��ҥ�wu����7-�e�QI���奮v��Cr�g���&�
9�����,���04��\wg�.����S��|b�C[.w@A�e?�_�ir�Il�~R���)"!�uްx�(?+�H3n��U�f��=�oE-�'�;���!�:u5��(ܹ	ǉ8X����oW�B�! >~��������H� ��5������;U��#�K��g�vd��H�A�a9�#��y[q���@��S�?F���׈�u7����t�Wݟe='lQ0e

�JWi�5�D�����Ĥ~E"�!sXlxVHYEB    9c12     df0�)
Kvv�S�"���y�)z��Y�E�gӾ0)��_�%�Z�@�B����D��&g�I B0�&��ayG�R���٧�BrB�h���%
w[�zD�&;dGo��_�kC޿��Q�?@���K��Mv��ANy���f�_.��m?-��b<�N�bS��ԇY�	���F����B3�@C��^[���F�ȴ�	&Qf*����^h�˷,��i�EsM�F�kBf &b��xF%E�֛�]"�`X�M,JV�0���Kh{p�mP�S%y�j���G����ݦmݏ��?l��|&�N���И�L�C����-�u�ޢ!$�,1�t��d��~�vړy�u�3El�ρ9�� ���as��+N`�G���<�m)<}*�~%,�cI�W��eI�σ��G�zܨ�^"�z��3� uvؓ�,6j KNNC^͛����2a����Ԭ)�
��pbV�,X�j�"u}AlGW|}�`q%��#�H˵�ab�V�GIEY�$�������tT`��7�c�T�A�6�+��<]�dR�j��gY(��s��-��"_*	�N�V�	�i�Ȳz��G^�/��[���2�+�T��Q�ŵ��h�J]�>3�y,ᆀNPO�jl���7jL]�L12w�=�����&�R���xO��#�ȅJj�y��N��e��o���a5 �[�D��uũ�CB�����&9񔓩�%3�~x�!�5���H��y
j͖���� �jv��a=J�AVHB�S��_�ܜS�ݡ�����e�P�3,
�� �8-)��8}sٙm�]�r�Wv��揷d��b�����KqDc9����=P&�+v��ѹ�v(�%^*m2kX�`�I����i�fF׮�M�����F����3���,�/fH�AjF�"4�s�����1e�
c�W�O؂.�^��
~L!�M��"��T�҅�L�h]�e[_�V�wF�~oN	��C"; AjCBɪk)��%�[��{B7�x��Mv�����\���*q��{2�R�Nտ�R����* ���\�b�n1N���ȓ@8l�.��e���
��R`˻.�r`�A�"PM9n�����-y/ɰ��8:�%��zV���B �7� L���F�N�<�׭�L�} !�]�=�k�݈�q065vñS�<��t%��"ɤ�"�{�ٱv��Sk!T�G�D��x�eY. f|^R+o�;�vȍ�����Nc7?�oe���k�!�0 �%$d�_b�� � ��G9+�X��1�?�x��i��F��~0�l첿�i��l�������8�2���'�aݫ�=�����*f��r�ϛ)"��ng��kUT���/-[���!|&I�"q1Gvt<#"����A�@k�{͊e�U����9�f�^��a��&],2�㣞���}��~z;Fy��欨�BY���<�|��ʄ
���^[&���$�:>�Z	!˸���|��;3$#��/ƃ�vb�r�)@�L#65=H���Fj�c���fɞU�TYh�9�DT�N�QT��ۀ�"C�Z3o�����H�L��P�8͝G<�V��i����=���ڛ�aWzꖄ�f�|p��0���\�ñ���;��41d\$�g��"��i��B|�
�۶�	`�3+6H�N�\�ui��Xdi��O�����Bʞ��W�p���?{&�w�b3�p���2�_ꁾ���*���_�5>u�'8��@�Oҫr�
E����������|#��$���3V�"Dfz	�!}�`��t4,�I+��`���*����X?C)�"*a��YT��%��3��� <4'��7�}��o��9����W�o��krƇ��;B���M*@؆ �][h(nAf��>;k�ϐ׺�O�ֽ�߬qi�5�`4 N�ά����#M� ����Ծ�0�����~�ی��w���B3:���E����if4S1���9� F�*.�Q���/����cP4gX��"�N4Ӓ�_`5@+����%:���,��#���*�y��ۨfzG�N�T?Up���J�9nV��[تÍ���7����ޞ��2&^�$�yu@c���kQ[��0@MB�	zv�B���)�� `+��`��rmhq�l�nJ�;��#���\1�9Fҗ����p���	�@-|��@A۷�8�P����Q.���6	J=��q��Y\=Hώ�`p��[�_��G<-2��I�f���zKSx�Ya�"��Fu��"?'|v�tC׊���:'��Oz>[�|�ȯ���Ҙ}��/5��A���^�;ݏ}C��ٛ����d�N]~��Wx!N�iד��;i�UL�'�0�:��Z��ê�}�����Z>_vz��|W3�Df�;���#���(K-���&��'������\�Q���|l/��#���O(�%P��ͼ���D!�	
))\��_�4	8H�;d]��G��;v|�Ar���>Mo���'-��b�m�N|���7�_�4@]1�m�n�mz�qH��dP�4%�-�������v�h\�ƭvC��dN��nj�+9#������c�.ڬ޺k�X
-Ғ��i'U��;P�����e�������5l���։`��E;B7C�b�!����)B�֋+��9����k+�񋵔�ce�\X�����a.��g|�Eȫ%��X�%��G���c.���̅�/�+0���m�l�!��!�{�:C�M�ltH��.@�,�vdyUA5��Fm��dl�^LȒud_:�FH��!� v4��f�@
���SG��C�߈(��^���G�tv�~�&�v6����P\��_{+�e��+ � :���i4���6b�7�e���ڈz~���i�VK��M@���&

�朳�Ŭ�N%͓��X�/��$���q��r�M��?ۇ��x�����r�5�*{x:e!&�Z��N[���C������3��~���oS\��UQ�'"���P�:"�A�������y#�$�x�X��B��j�@�g�$U�c�[�_!)��^�]����i��Ev[ckC�|�)�q#1J��|�1"�wꒄ"� q�_vRNH��A��h��P����ֶ'����%����4��I;DˁQ���+"tT�D��r,V1{���QN���=W� �_��t<�V�E��:lAz=W ur�?7U�oʚ�I��Py��/�(�ǿpe���C�2/�Οn�ּA��������?���Y����c�c��zrbO[_
����?:����N| ��^J�X=3�2���Fp�G�������ζ+�O��\y����ƒg�͇�B<e�{0mV7����T�v�q	���MH���բ So���Z/t!u�|����<x�c��*�*�_8�rV��S��Y+����UR����k >F��\~�I�ÐF�oYa���z����"T+�ܜ�6VX��7G)��h����50� 9�,Z�7�qwMn��V�=�C�J��e�A�&���_��/lR�Ӈ�%����D�