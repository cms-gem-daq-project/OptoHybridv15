XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��uf��)�M#�(��N� �!��k�Yj�u,0�HG^�eN��6S^�K��������ł�hI.���e�z	� f9�T-�$�����0/!q����f��|���OM�v:
ـ�ʄ��C<csW���-���
(���t_`le�_+h�kK���e��1T|�N{\ƞ��h�8��ϴi�w_6���H��i���^��[������Sƺ�����Q����+2�(ѽ����UfK��e;�3�Y~ ��
�L_v���!�\�2��W�g����-
�k`�n���s��1���3X�n"/�JXO�nJ�.aDl�+���-Ьu�����Ạ�u�t�&�Ȅ�rg1���Q��e�C����T������<ȡ��L�p�ͱ�����"�P@j���4�~�������87��&q���a���/V���p��C�;í�%S�G����X���]��#�RV�Nr܌���"�C���*߄���Z/�N�qt���=��.V���}\L�0�����m��6ά
����ā�!)�ó�{ F*4�{/��ͥA�cX1̠��)[������I��ۤ���'�dH�F�h�W�#7�q�S���\���k����=j��$��N��a��-'VJ���r9�ݭޗ���W�x2���6�+��$5�4�P�7lJ@������1"�i�q�ڸ3Uu�r?�����G��zia���Kc�����D��\�Sf�x���~`q��ߑZ�ma3o>XlxVHYEB     730     2e0�9j���.��Lt�'j��9��O�
�r��$^֮	��l������pXo���$D_��n&�?~sQ�`}�7�ċ�D>e�[F��N7�/[����>�cX%��g��t'�'[��0�k��;��
��s����?�{Ꟁ�%�����S�>8s���䁔v���␊�%~_�ken X-�p�����ޚK�nqӚ!���,�K爨Ҥy̽�^Wl���f%��M�hNx���[P3m	��۔̇��4���$��BC�1ǐ_ �8B�D��$~��/G:H`F8G]�Mo]	=�=v�ƽ[ "[s�cZ���6E��;���+�A��7�X����Kyfi���Ő��T*�(>����G,�P,�
��OqS����n�I�&��f9�Z��ݕ�v�-�v0�l����mijU5�&������̥�=��}��0�4c��[�5= ��%���C\����$�9@������3�n�;��.��HPdZ3p@D������l�1D(�=s��Ds�x�(�Aus�p6#��?������l���`}�E�ѽ C�
�<e� ����}z���I���h��@������Fvؐd���U�+J��,G�k��
�m���-������/o'�� �xCh�%Y���������,2ґ�����H��l;f������Ho�B�j�!+���{G��VCSd�5�(��