XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Al0C�ֈ罧���b�бA��f~�C�F`#"֭Y����c6��tdA�݊�����)+SL}YZŲ��~y��m�Ożx&��}4��b;x	�@�dO����$����#ߒZث�i�(W���1�d���*�h���-@�����e���*���L�y	m��&��y5��:f�z#Iw �*!S~k�W�#�l
�e�N'�O �$�vpƅ�o�6u��C�����3�8i��i��\Xܷ���O>�P`3�4^� ����R�i'z�-��b�4O�_R��hO�>�/���EI#�T7����,��E�9tO�tO��'�@�z�ҧ����D^n��&���h-0�L�B�0{J��u���
։�|�>���E>��Q�Vknءj̴"¬l���A{������[���(4�k먳b�-�V�@�Z��PA���>�^��K7&�t7C�Sku���6'p@P���U$�)o�!E�`oмm}8=�n�2���o�߮�fj�i�Q(b�2O�<
J0T2d����͒ l
ނQ��J"��BT��O�9��g�� �ժ��u�����Iuhɖ�?'�ŝn�@v��������IN�[׺�F�J�-'�RQk��Y�"?z���O@x�&�+ ��Z/AV~�r�T��l��ů�?�=%hv��D[��SW�6�s��%Vh�X�!�Q."�o�=��f��_62�u$�=*ŧ��Ui*��'�XlxVHYEB    1c48     560J��¼ʪʝ�r|0�S#����*���o�`^���`�e5�	ϔȀ�e!��t���0�Aۮ��ٛ�9k�{���N�
��M٪a�����5� r(¶��W|0]��`���D�� �G��t��1�Ɍ��/��j��B��¢���E����׿�AP��Z�1b��	y�'�;8n�Y�xg��9�Q�묂cq��L�m�v���2��'��7l^IFz��*��N|�|�-�>�v�L��%
�O;Ij�-�\�<Rz��R�g�����I|g�6ޠKX���F���`���K���I���#�z�A��-��4H*w���;~p�  q>�Z����ۤ����t	���k�Q��<�h�o���\��ԛF�	� &�`>���l;_+��$�qn�u�{C�7s�,*hԪ�l�|��-Κxo�
no;%�8�P1˶rT�è��k%6S:{�'�p<g�!R��JE���W�����(���(�44�V���К�9W"w<��L"��o����򝴱[��l�/[�Зe�:�3{�����{��?�3<v�~�x�V�J�y���[�g�\���Yv��?Ċs)�r��M�~���]h�q�K?�.�ؾ�ȥ!z'��P`�t�����Q�����ew�����!��;��â,�a������]��������-\e�F���Ϙ�A�l�*~)i�0�Q���a�՟r����T_bL������;�% �9�C��#P�w��F����y5�&�����ب�K�M�Ւ.�fg�K���Ve!�NMe������rR(V�
k�h����d��V`s����}�A�[b�"J�Wg������7�#�4,�Z g�y��[�]��S(�kE�:��#�~F�Tt
��ζ\���#���۪���/5�ˮ�3�*���lԋ:����7��#^��z��-���� '�,�B�Vw��r�X{0(ꟈDth�=�K}.�7�L7)r^iq�2�h�#����4S8�wLN���+̄����{!͊�I�%�����-�\Z$���yNiV(-j38��}�3pV���/�ȭ���-8Э9���"�g���ί�8m���m<����Y	�'��r;�:�F
I�ddtq�(��jl����۽k�]c4+J����?�Mi1����C�M�VD��Y΋��2:���##���Re���c�Ac?��5P�/ȷ7C��+pJ<�� �8q$�(pu/�)�|�m7F�ƛ��M�0��c66%P��$��a��1��5�s����f9�#�[�s�Y_a����\��Nٞ'���p���5��x+H
"ND��SKj��}k#9�8������