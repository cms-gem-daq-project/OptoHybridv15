XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2�πk�ű��s
gC˓�g���.�"2y�A�Z�ZW�L����1R��̅�B�_{3���|�fh�a��$8h�5���<`||�g.�Z�`$S�X8n�
_�_�d(���8�@۪E�>A|����9���6D�%�6�����Z;[��I������ľ﮶B��Rn�1+�f;u� ���Z䠤�����!�R�k��6X��0��+�bk��b���i�ݛS��K�����`�LV�n�� I]������.+2/k.DJ�c�]U���fe�s��]�S:���~����`��e*���ᘠ�$@Jp����e�#�36�N��{�LݭK�fn�O�.�"�!�5YO�C�u��������ȇ��Zx����/9.�VQe��2����3F�`�;���6�� HR^���a�uك ��Jh� L�[��;�����ۅq#�ҴY�B�}o`
�*5<��#p;)R�� _�e����z��<��U�.a{�8Z��
*�a���"%g�	H:�s�W�?0�$��a��J�Y�6���q� <�����h�5j_�88L\��Zt��mٱ�$�nS�����$����$�Xa� J0�2�nRC�C�q�J����ˢH�
o �є�f?#�tVp-s����$0E��zX���m �}0:ow@�H�?�>���J�j��RL�l.d �i����9����zd�[f%8A���H�ݔ[�c:�ßrԍ��S�+b (���!p���fXlxVHYEB    690c     b10ō��r?1�{2\�jm�B����b�Xn�o����y+����og(�R\���u�w���(���ɕ����GtYXK�S��s��1$eW*�<矄�,?5�A3��ۆnܵ�[*e2���?�6<ˮ�w�����;׋����je8h0���<W[�i�]m^�{�WI�0���h��]����� ��N���樋x1���9�����xx�!�(-��
0��W������r��)��v�es��e5�e.��;;���P"�!1i�W�~��{EZ�4�Ĳ�tT�j�')����]�C(�#e7��`v=�M��YU,��3.�\�P�+_�7��P���(P��i����l�`P.���T�H�J��X�n�/�����f0��g�ړ��٦k(�] ׸�s9h�f%��E��|��f䑔D��:np3�`��8w�rɅ~����#5{��(�� ��xT�k ��/��J]�:��b�)�C2YS��ʵ�3�jv�bQ$�^\T���{��&�~S�~�O�Q��F�S���7YB�a�,1{�[��ߣ�-����f7 2"6<�4h�t3�\~Nzl";�������;Յ�e&���o����Yꌏ�ÄЃ&�/��ب�;5:48���o�����'/��A
�V��s��-e
��\U�l�����t�o6�-M�Kx���2,�φ��	�+�Z³��(����C����^��H(��EV��O������%�4��Y&v�nWtSY��8��w�a�����ц�)��G��,����;cKV}|�pf���9�� �����Ȧ�5i m�W��}V��3���\��y�,P3�~�	� �s�F� ���q���If�+�aS?��b/�v1�ȜYA�B�`���=���0̙)'�n����&۞+�d�=2V,I��D�/������Gό҂���Զ�E���lW<_Sb���N�� ]F#�6�#[��i�Vq� ��T������t.�T���B�D�D{^�y��n-}3细ʥ��IVG����EI�/�5u�������
Q�uN�{F2�sb�99A9?4��9�g�^?u��l��@fG��XJ�"��Y=&$��Zu#\�L0��E��R���z8Q-��	��\�r��c�Tʫڎy썱o���S,�
vl��g"g��lӘ ����֟ǋk&��X�8�!|�3e�o�ܑqM�T����!l��W��[�8}�s��4k@�/�>.%����7F,va��y�f��M6l��ks
�o���˱��NPqu�:�  ������\�2|�l�$!x�d߯�ߣ$�2	�_�����LJ[��>�ծ(��B�*E�&�Z�Z�(���Tt�02B�+�bH#�g��ܗ�FӾE!6n��*F�oN~^R:��d��� �8�T(ԡ�������p��|R�\s��0�p���
�u,����L8=��q
����2i!ӥ�U`t06�m��m3�k���X�?&�
�`I���f����&��RQ�B��bu�Y��P���ۦ��:��3�%�\�]����	�ޫ�Đ�=,h2)�rXY~�܋�,a3�O^�6�U~��߿z)x$O��g��;�9��M<���#�zqw�	��Df|\��H�R���Ն��Qn��H���Z9�d��٬���tQ(�P	�s�-RU^��{Br1�͖���+T&���-5?�솮P�AD+����t��y9	P��}��~hnտ�����Q������-o�������s��WZ�F��\��?�E�ҩ������8`��lҪ�W�ܿ�Ļt��_��&=Bgޥb��������<�6� ��*�݈u6�|���o�z��G��7�����i��*�5���V� ��z-%uG��,�CA�;��h�H)/���Mep-�R���nQ�4�N6�5��(9���O�6ɕ��3LR������N�n~c)B�RyH�ĺN%�}�	����;��
 5�v��A1mwx��fܓȺ���6����tw*}"��hL��T�
3�Myܴ���,��~O��g=�9n��Sm��a'��&h9���sR8o6#��tX��oґ��Uҡ�O{���J�� �m�4HI\�:��mV~ݦ�����MkB5	Κ�%�O~`��8\�n'�;!R����t#Jn��Mi8�.g�(��gI> �Ԛ��6ޚ��M
�U>5+꥞�����Pa��\�4���ߖ ?m�ӊ�ZB5���.iL��nj�/w[~�S��$J�7�x����b!N3ڡ�X'�J��!r�\�s�H�,�g2sY#��:��j��UY�g��H��y֐�Ȍ���ZP�%3�a�!�>��v_6d��V�ў����<�H���������
��ӗ�
}����!ֱv��V�������L[�j��g��K�c��z6O��V�4v޾���#�K�B-O�E�e�6��^[bJv m5J}���$!â���:}�����w��F���b�곿_�X����\s�t��2��1YiHn8PC�J��ؾ%���*]4pz�<?�D[���v.60�
�F�8^MX1W��V�;�ú��˭�5�橄ʫ볆��8l^#������d|D�,*�"�H�/�z�煛�;}	����;v�b�^�8��98UX�B>��C���L�A]Gꑇv�!C�_|�@d��1߼jRw,1P�Tw��ՁVH-C�1�ƨ�C�Z�Y��jd�Ȯe�TdL[�0W)'�:��X�%h�