XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����u�*ۆvEV��k��R�廷�⃚9��L؟lٲ!���:�B������߬{������O�P�t<Տ�[���i�x�ٗ��.�
R�f
�pmx�A��ܠ��b]T�~���!Q�Ҫ�BP��Y��7��,C�D����;��Je��jٙ�����<#�&�lp�[��Ԫt��=vF�v�p+�h7�-}4����3M���[�}ٜ&.�6�f9P��KR�r�r�H�LT�̶��6M��5����7���1o�	9ki[��K��6r�7r��Ų71r����녌[��H�O�h���:��"��ͼVIΨ���Qק�&W�Mr��@��X�T��B'�<$cz��\�+����᝹jc
&^�e��'����&�������F�֟J�M?�|�w�)���P!ǧ(���7c�&�7��]�2���S W�ֹz��Μ�m�������O��;�f��.�U_TeI�Q����z��?��6��b�S��F6�c\��ρ7��@{0bė><l݃�G$l��aJD݅l���0m��Q�%�Q؛�v��Ϭ�3i^#��u����S����f#�Y�4�щ$���vU#���ԛ �i`�M�}�~c�^E��`��k�Qg���A�9��82	�|1K��R��z�Y=����D�>;]�� �F4��/}_y~|�V���c��a�>����
G�=���p*��[�� &�����yNuPԳN�mj���MXlxVHYEB    1cf5     790��[�n]��!.��#�B�U���HމYp�'�u߰�i�e�I�+�doL���D<�>����*?�$x���x
e����?D��s�4���:�U��w@��L�Ad��ؿ��IN$��;���p�����rņI]�G��P�v��
��~�SD�1X{tc: ա�!�OR��
ǜv]gdV��a���`j	XTE�dF�j���Y�)�+ ��0�y�ړ@�
�Y�	��d��0G�J0�Cj�O�+�1�DG�a
�PȐ�b� p����1qe��n��9�s������}�V�Ҹ>Ó�<�0��[���2P{�i�kv�h;z��w^Ґ��(���ws���<g��C_m��'�8����ҡ�y���'��T�����>V��f�˅�;�_5��5�1��'Mk��S=P�n���Q|83�j �=��^���1��P?�;h�~l�oř���PUAPi}����G�!4��G'��ܮ�A	�Ṽ�xik;���^�ܙ�>~.B���H"Gm��9+,��mR#��|���b|���2��� �	v2�r:i�U��:7�d#�bEl]�覟ĺ|����I��ԭp\��X��,\��b�TX��!&ɕ[D�?L�G{�=p�/� �� K���K]�G��-�M5-���x��� ��A��VQ��L��Y̵fY��_�$F���v{���5R�{��)a��\k�^�H??�kb�XH�ج�9�~g>�s]FgU2 �x!B�]�+oء�U/�G��G	���/�(XZ.�a�V ���w/��D�\��^��/htiA1&C� ~�Dm�K"�R����,\O�3��� �FeT]m�"���*@��m���3 ~�5I[X]ڠ١���K�gV��� r�>-�М��6�#���*͇.�N�<���2��cl. u���Y8T��w 8)��W�[Z^ӊL��42����V�'�U�D��4�u:6C���g,��._�aA�f�#j�����\�Wj�����	*����)��h�s�A��5� ����1������$���a�iݦ�*�� ����gR���؞SRw�YA�Zg����xzf��D�D�>WB"l%���-0���>��PӒݡP.C`�L��-G\�v������/�b�z}�.Z�o�wۤU���N�u4��Ⱦj"n���e��7*C;e
��A�]���ĝґY��+B`K��o0�8����xB�ڋMRF��A՛��)F=|蹔E��E�k<%�7A7�ah������&]���k�8���O���8���4҉��2ȡJL���3&b���J�r[��5��w�.�B���a��J��`Im�tZ�� �,����B���LY��	Y��L1U�iI�����t�Q�Ƕ2��ʙ�q]J�"�ȗe��w��*�CYEє�cS�?b�@�P�|w㹵<wi�#īw��1)�w��N+ P��cU�e\��ú�?.j1P	׽��&�~�+x��e��1Liז�KM�	�J����=��Z������]��R�!��2n�T,��ˆ4C��T�٬���w�E=c�p8Yr6�45��CxzS�~�,�$������A�"礍U�^8Ί3f���[�_��XG��:�<��^���.`�4I|����q�9��	�tf�zsZܡ����;`MX�	/���@i�_�L���Q2K������q��?��s8�on��gK��ݍ�O�2	tO�$:��c+z�e��<�������ĳ�����ڋ�-�ò^��ǩ��F%�"ia���8]�]�1�=���a6�����Q,J�"zx�o�~�g�8�5W�X��=�`ɀ�&0ZDldp��ۍ��A�����,�[kt��&���Z�{E��ݩ���9���h~M