XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��QP���	|��h��N˭�C,Y�uP�>Z�w�YH�0�證�˅��;,�F����9�XVE��V��פ���J�z�슪Ճ��x�bR���Y>�)��&B7�0�P�\;u�"ݷ&,�����I>`�s�4*��c��"^'˻U�3��Bم`���bt�Ɖ��w��)��vhF�BÞ �����7؂b��'e ���y��� d�O��(���7͟~_��D�T<b~Ԕ?7*�ga;�qL�����+aEc+LO0���M���O6��+�tB�_Zc2�8k��)�tC�|��Dn'�3��Dix���z�Щ�J�#�]z��ŕ
�4�2���D@3�+'�m��T����`�"�]��D!=
=���Js�����9�C� ���ԫw��&�
'X�2iy�~�ni�C�+ʿg
4sO	��"�x��>K��SѢE�k�>3(�g��3˔���hV����He����(x5g&(����\�>ze��ޫ|��wp S�$AFO����{�C������C�4;�3rT�i�"]��b%7y>۲���^�x�����P���PF���ZD���;~js�W�{���OI{a��T@��.��l����6ZY�-�P8l2�t}���Z�B�V�Y( �FA*�ڨ�����x7Z̪���즤%cHͧ+J'*��Iρ��$�L�ta��\�0�S���JN�iїT �AI�	�t�}S[��CVp	e8�A;�W���by]̷3���XlxVHYEB    2864     8d0h T 0����ύ��*�)X��d@�q{&<����0�:��L�m�0@�����Y
F;��7?����N\L�ĝ�ީ^���#��8D��P 1� �?�3�pӖ��}�2�2IO4�{���趕��/wk�U#�8��_5���dY;8��?HH���9���_�N�]XP��𘞤سL�9�s
D��Y�F�p���0�ʉ��Ee�������u��4�Mq[�3��,U�
kJ��=&�.F�/a����5�
��q\7j�}���`0F_����~�<)�)m7/�y���\�J��+��Ɓ�K��VƜ_D4׫���uDb���4<m5���W��j>��n,ӟE��k#ׯ�>����Nko���٫ܧ��_�ٹsg��F�P5�PNct�vO���C��\��X�>+�Y�&�o0N�bA�0�&��9�r8Trh��qX��fLʒ�?����T&k�s���K�b��8خ�q��}@��;�w�?3r��-bT)�?fgZ��g]���UH2���K|G�L�~(����̦�<�;������Wew+Ith䰎;Y�<��Wׯ;�ҡ��{���_�z���f$M9��t����u\�T��t��X&��:�A�"}�J ��-���D����[��,�!8:��o�����磬�|ϔ��j�::*9gLٲp�x�g$�.R�%"��A���q!�kw1�5<sS�c�&���"�mnB~<yn_�Қ$�6����~A��u]���a]��q�x��-�bc�Y����J�㽈Z{�<�� ���qt����E��^�#=J�v9�
�@�"����B|�;lB#u߿����W���47I�/���(N����Ǧ�ˣ唖K���1�	*�c�8�h�i<G�<��k62�m�����1��P7oI��*~�w	�Y�msg]Cuo����dY�'�Z��Z�騮X'Q��%r�W���T��l]�<H�+*WDe�\�	��$��ɤ��E��-sqJ�H��Z��;J��BB�k��l��S+�~��;%z���enjQ�*�%������c"���e�o��[�"�8]�Ǆ��]8�d�v��Cc�9�-x�����B���x��m� ����ӊ��׬��9�țZ��sA/zr����$�T�6b��t�᷶�4lcT�=}s�
W��!�ݣ7�5��5���d[H�j`X$���4�VY�'=q���nS"���"4��g6�ɸ�h��|J:������g;�t*���G�7�mɨ��x��5�7e�U",���K���Rp/��@�3�IGw��)�$3X������k�P���' �ٷ��J���(Z�]��jm��:�Zֶ��Y@�T����'. ��b���{	���kꀃcr�I�����g=Ȟ�
ʻ-I̧Q�o�>������vTpz��IGZ*�8�>|qj���7��|-}����@��a����a2����l �-&�/"t�"��e�Q��nc�V^��j����͝��������w�7��ؐ�k�'[�s;���d'We�:\�����G�5�ɞr	k_ByE�;\���6ԑ �z[�ƃSܵ!�f~Vh,�#y�g�6� �Ȝ���m0�K<~9l�J���;�4�����<	�J�8v���_�UY-rRN���ڔ_� ��oG�[sW�C�+}��q��8�
6Hx�5��"��Sg���
�}�T"��ϗ8V[�]D�k���ؔ0�e���������$FȪ��x��:����B<���3�뜖����q l]��=�R����n����+ �@�2a�+�B6۩w��Ғ�`I� VtVB�N-`n	&��ԃ�v�r�į���,�l8�,P!a��)�'ߐM6�qV8��UD��U�8Q��eT7Uy���w�
,�)�0���#wV!q������AX���5��Ƭ�8V�[4�n��E�^4����S��[�r�Y�?�J^�>�1z�"%RZ�m R0�J+���
�1)U;5�_LV%�-aĆ�n)�_�F����U1m󰔻�Y�Zm7x{y�c�0.0��qB���#ȾLY:��˛��J����l�ǈU�c�dc+�Da��Q�o�TۯY����t)i�#S�오1e���!�A3#h�����nF�3OüZ�X��� KJ�(�␛�.ur�g/��*}�j���6j�,���n��m�=Q���/,��1Iܚ�8��8����WB�T���EFh5q�oI׎���,�|_&