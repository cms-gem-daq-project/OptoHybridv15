XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[4�	.	���#08!������o�7T�g�y���hy���R���ȯ�k��l}�Q$�*V�[SX��l�GC��6���e��_���:�M�Ip�V�!cU˾p�&����Rj��T$�O�����f#�-3��9/�KI^�"d�OW��BL��n�|}�h:�?����[�?�0��	����<�ۼ��ݸ`QM(�N��v���x-��Ta��}����	�&"ϕ��T.�����C�D�u�Z�Њf7���qh�hpZp[�Gy*PyT����^u����卿@6&���/�O�y8�����b�0;��[��!�S�.O�ʒ�~�S�$����b�d5����5�����+�۾��c6����ZC�Il&v�"\8dfʧ3�?oM��s=��FF��X��}>����C]t����n�"�8u�����1�ך$��N����I]�����	�4ЙT�O�g2�!mJz \#�źK�K�,o��O���
1^"�VH�cIbD78�f����ʻK?ۍ�X�t�a<?���2�A�4��zO͌K�aD9��	�Ѭ��1i�Dp�w��(�bx������A�҉<����#O`�t69��(K��^�9G��0��1B�ۖ��٦8���͈+/s�V�� ��w9�6��*�������>A�d'`��� ����d[��蘸�¿�?e�mx�+š
�}���kƝ�iA�Qh�x����Ձr�6�f���xD��������(#e��ĝ��5�_�w�Wl#WXlxVHYEB     7e5     330�����J6�Ҽa�3F�T�SD��Seq�-S6�Pre�>�]9�3��'�/c=y)��A���`���:�l��P���A�0��r#�9|+u���n��I�H��t\��+-�!��6>��_Y�2��0[���dW吤Cc�{Ǥ�ƍ��/�/��~�6D�~�m� ��:�'b����+�*��t.��9�d&��8Y�nVgQ��V*���S�@0�"�U?j�\��BpT]���%Cg�:C�S)�m֥H�W<2J�9�9�M�` �F�gWU�BQ�~qΡ�3��{r:���[����q��z�����'"؊���1q{=�y{d�Ó�?��è���B�+���N彉V�Λ�ƌ
[c���_=��������*ZPL0��" y�9��Mo��2d-�1��*���q�Yix*l�RA'�@~�WR���x��R��������72��98؅q4\N��(�|˽�P�f ��Ƅ����m���(Xڈ�eij�_��ʧ�_���l�U�~!�Ch��^�gt�b��`�c[
$zz���]l^'I.&��u�5�ns��e�U�8����R��M�ĳF7�]tJ]ޑ��j��ό�O���X���2l�i�<��w��·�����c���{w[��F���"�� �*�� ��hi��1�3�V!�q�����*�y�5B˪�/�!���Ё4N�W��S����(�^&�~OfC�l���'Wۜ�8p���9����ش�!?��T��OO��U@bL�H9K��F�?�3Y�~3�#{�mG��R��/�K�|{�uk�U�Y_�5�&5flg