XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+LpnwD�����|�+�5��i�Z�x� �!c�-�j��D;�+M����v�5o*mL��c6�d.����AR�������;*��Y��t�$���������X,�i�f^�������?�肚�owv=���7ճ%�B0BP�Xiq���W�Fn���F���K�u͞������b��5�,�NH-J�
�P.�L��4^OjN�4:���~۵`��aY�����;1�@�/.`A�P��@�#A��W��:���mxF����],�E�?۹��̚���|-ۤD���*�I)�/ٮ�g�0C�HR�$�M���@�Ôd��șI�㬣�Ƣ���H�_�$@����U-�$s<0ͭ���T�.����L��*����m~�����@�]�˶��<���aI�Z1��w<�D�+eyk]�����m�2�k��e�f,{�k��	l����fx'%��(��Yy�W�WSa��U�Yfh��j�9�vC�vo�4���	��!s~-T�y�f�1?�2�-z��M��e#�b�mօ�}f9�����f>Q�w��e�Z1\�0�'	'0Wh�C�`@��m����]���=��ց�~�����W�;�]C���.��'��D
U`,[�.6���:�wv��)��k��̡س^��I���[SZB`Hm�Z�*����t�qO�h[�s���.y��f$��;�+� %!��an6W�{�@B�}��^%�p�]a��u�3��VL���(�lK���7F��*���XlxVHYEB     686     2f00��o�c�� ��>�k�����rl�/�L���S�x(���F@��;���PR��\��0C�i`%���� ��.z��S����cM��B���D�*�0���]F+�u�cB6���3z�1�w-��"�@,�牨I�3D�,ס�R	�U�u����r�l�-x�O:U9-�k�8��!u���o}�gR�Xy���s7��~������ԩ"�-�"�T���2�ZE��f�N����>���+�p�������@-����[�zfʼŮ�g���mȀ]E�v<8�S;F}�WF!�o�r�pX����`%�� 죞?#72Ĩ�#> �=Y�w��#&��F�D���FG��i�V�QV���g�/U�0n�LkG���ܶ4�g��Y�pqɚ׏�I�;�q�����W�w��M$�J���rI��+H5	%��GĶvIw.D���@J<��;i��'�S�_��$�3�g��O��ñv��?���d+ୄvqQRr�,U֓��S� j�̞�m��e ؎i�j9�A����T�d��Gk�ɨJ:NcV�:�������v�O���Ϳ֙k;$'����+%E�p|5S*�3�����i�ͤU�R�U��V�8�&{�r�R��<���G8��.ȗ%3�X�Υ�����s�6���.F�������`ע�����ob�2g�+��|^�0�T��8^A�� Ѹ<1Beb�N��* .��)!����������W�T��+���ˣ��<�\P���;��C���g