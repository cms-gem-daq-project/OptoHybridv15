XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&��>�D
����˾h0��a�����kt�������ؚ�+#Qah���	���p�����0F�����޴\A* 	jr�y�ج_8w�D��o1G��ϚTy��*�	�M仭��d���u����%r觡ꍡB������i9ҊGkڈ��4�g�uA)D��uo��[�Q������Î���6�;�
nk�'$��s�_�!�~7">��������ᡷ�+����P����r��zj5�~�M�
���{Ӡ)x*�lk�����B�ɠI�<C}/Z� =�cSfAÆP �o�0���[�k3g~XuW~�\Z:_CO�p}���1#�h�A-6=n�;��7�&���<����	�&�9���Q@dh-Qc܅��>�ʿ0�x��d� z�(��Zi�������{[���%�0��cԳ(K��tE7e���t���� ˲���w�?���[���m���K��_�P�z��Ͷ��&:��!�ed�m[/�#A玤���r$D�Ƹ^�'�M���:�r��+�.-�uBK#�9T5ܺ�}�@>��؈(1��C�H3Q�bt$1T��^n�E�Gl�|�HfR����os�#���:��Nb)\��X:�u	�G<՟˦�IN��@��jw����ǆx�~P �܎��GU�q0�-1�b�{��A1�٪�l�zH'9�a˛{��P|�MȐ�wZ�t��;i�ԁw�X��_h���h��GI�oC�,%�����1��#��������]��"��tN��{y&XlxVHYEB    6fd8     c30]��=9;UP ^i+���UG��� ?R���<ު�<]�M��J�u�u��χ�"�\P,���V}�s�$�-db�!�HK(k�\�O�mV�, &�����>(;Y��Ve��F�JϾ���D�y�,���N*$�����2"H��gC	$�����������b�~=�\>9�=�R��U̟}A6��h�k��k���G]��׾��2����������N+�(�#
�~5��Cw��0{��LP��Q�~$���m#3fqz3zPcϏ�"��]��T~ z{�<�ϥ��_M��>�5����m���z1KM<f��`e�n�a�M2[ǘ�^r���y����	�ݻ2(Y���%d����1��I;�YRR��<$h#x����;|5TKO4e>7ϣ�����dwͩq�.㩆��O�����+�fTgc�dBm�F(��+��1���nE�h:��Ws���`?�A�$� �fˁ���<���5J���z_�b�#�~�AԌdmXuU˾�;t��A�x�l�N�20�B�L�͇5�0`�}���m`֚T�;��qju��w,�F�0)�Z���?+W}�{q��h�����c���.����g�cE�&�F�������L�a�Sߗ��/�+�fϓ���ރd"?��N`��g���!m�����B����yÕ7w�i#w�
Ʌ��J��0.E
I�y=M_	-q�:�P,��{�}�~�h�X�0g�����6�)�n�L.�o����]zf{b0c�;9�F�nIƲ8�\��$��a�*4�Ede6�r��O|��T,*�Ԧ&owFi>hp8����wǴ�ъӤF~�y�?#yY�j¤��9���B�l�
�t�^Gqu�X�X�O�S��\��������V��Ms��9. |2kQ����OF���H,�R�tc�������a9��4��J͛B��t�G�"�^��k�������X����WN��g|Dۢ��2���,��!& �Ɨ�b�]��S����4�ɟ��3��E$������?�!�<(�S�\F��1ir�/���i|6};绉<�ʩnc�IO�&�ht6[N�'��al8V��j��M�����^��i㟁VGv^!���\}I�j1�-X�{U�=�yz�Wp�:�Mz�Yr+�te�g�(�;� *���Vk������fv�oτي�4%��o����S�[Ń1-�y�E�Rl��'���J�9�.���9f(l E�X��f���F��L�و\���,l��@pc�1ᩣ���������l.P ��Y�>�Y�#����N1MG�k�vW7��q��ͼ.�Rֺ-c���7��Q/��]��F�$c{c�;�c3I�{��>4�`fM�Z�|G]0m?zH`b(���]N�k"�=qo]���y��X�# �+\�Ɖ�6 ��9�Q�4jE�ֻ&5yû-l�=����3Z�=̴b�#�	:��e0�A�	�; S�<1�&���R1?�����i�J�� b41�aJ5��9������[�tzUy�
�o�!�t���p,��4o����� )�W7Ƨ����-|Q=a.�E+E@t�fiO��e���'�zC�E�Ù��W%�P�\��EA?���}Kr�i3P׎�HUҵ�bȆ�I�苃��)'�Fi��u���G̽���B�낒`�y
se�h��6���~P�cxH(s�ݨr;�{-�����7������!W����YU*���d�Rkrd�	���P���Ҳn2|�+�|/r$�
�eo3�pJ/j3o�[n�������8��{�~���tv������"^�6�ﭟ���U��<�+�|&8iP�r����E}"z?����`c� 6O���2[L�C�T��d��Zit��%��UM��fF3e9;�����W��Sj�R ?�I&�������RX9+=���������mk?lU�o� i���|�NKu���btEA�"�8#P�9S�HF$G��׆��M�r��|�(�X��1\��Wͻ�ք�����͎�^�AF*���VA��=.��;O�����!����_�h��^�/oBm����h��;�@C(-�����;9�Q��J���A:���]U̄��Pw�#־ea���H|��H)٘X���� ���s𪻳e�&�'�h߽h�_~�Z�N�qq=�4O�g~�L������œ�559�F=�ٌ+c���Z]=�\����ɲ׌��]kshĬ���¸1�}!�X��_���<�]��Vӝ2
�#��b�Y�#�3�)f��<���8�z����eq5Y���H!+v%���#�R��byԯ@i-��5�s~�t�@lƵ�\��~Lv�*�N�eU��e�~�����W�.�d���,9[���
��MF*���(��C6b��T<u*T��渝��IQ�%��\�\y��W���*�B-�ed�8 /��eI��.^Y�p�����1�B*U'��R.��Ӆ�{k�̿R�k���c{E�����.kBbP��7s��G�T�*��/�ؚ�/�R�{6]�UVЫ��.�H���� �A$����P%�`���BKD��h��A���UA��Fg��sE�\K��C��|�������/d+�K��b�e(��O,��H�3�m��8)z��a��X/�#�Rm�'ե��?��+�/y�0�<�����Y9 Z܆��^���U�5�7���xN��X� ��o�q0o�� ��3w��L�E���b#�57�EY�7b�I��P�S�m��AY�Hrw�$- �(��a������_[��@,.��I<\*i���K���qPf*oU�F#U�>���Luu�ơ�lϷ[L���b,�~�&4Q�40	�X$mH��r5'�RXt	�$�'c�E���y��f�1Q�^�<�m�u��*��>�B�4I�!}BŐo<,�i��=M���+����nAl&s�=�Qw�4��l(HgJ�帹h���d S��,L�4�!���#0��	Xu�{O�?6>��E�[:�}>�g�+L�e�.�|�ɂ�𨢴o�q�����d"H��Z���7�g��Im�=�