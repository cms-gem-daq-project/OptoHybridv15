XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(n��2��P� ފ24 [p=�C�&�xɬ�S��&��p{>L)ِK5�^r�E����x�r�Նu�_�!���Khr(w���-85��3�y�m�0�,RS���EeN����|�I��՗����zTF��oȺ`�0�����X�M�@�}�r�Í�F���E*?aM#�XoBi֝�~I�ECs�T��?~�J�\C��K[E�Ġ�tU�a���sX�͠-AΟe��� �[)�9ڛ`��&���yhm������,D����_���ւ�]?��ޱZ�	ˮx��%��ك���G�Խj��B�0=�6�ŖO��T��;7�+�xE��B�ګ:����x��Z�@� s}b�~����Y_9w�$��m������|�QM��Oi��Qg[�V1�B�5W����5 [���"J�|Y��;5t���ٲ*��
)�7�qRV�Ex�C��Ń���E�Y´���-�[2�.4II�S��Oȇ�5�����5Q��s���J�����N��X����I��4޼�ϖn'^4�q��3B�}H�t
�<�r�������Fa��*&������$�O� ��Q0��T�G6
QDhI�^�e�rf����gh�]��S�Ȉ��z�~�b������� ���ձP�6;�5ϊI�b����c�=	��/�{��	�<s�
��}�dǈ=S���J��X�s��� �`�jn�1鸛*b��O��,����֍���פ�~�H��LH!XlxVHYEB     b08     3c0������Oe D���8�#���HVb��X���OJ�M���ܧ%��
���¼,?!Ա�'��3^�_�X�6��r��v]e�4��;5I�p���/��昣�l�2��P]�N�=E.���C�:	�,�;�!����K�{k���*���b�E{�j�S%TB+^o+�-9q�L�{�M�Z� F�{c�|��\��y�ܲD޿J����n�O�f�bK��(^{
�v<%j����e��ѵ�⾐��[���?���c�d;�R����Kڎ�g_�D�\O[|�8��}�q�� i2s2�l!��I_�U/'mO�O2s����=I7��4����Y�N��g�_wI��M&�fj/�� A�>���(-�I�d�{g%6��˸��'q��r�̛��"֧��K�Z�	���S�:��Z�$b;wƔ�S�fZc�����F,%w�O&��T�Tl��W���7@cbd5����#b�i��2�	 ,q�����[�>�<��؉b~4��>��b��1N��b_:O�4�Ƒ�����\�M�hr�L���D̬XP]`��k������ݮ0��O�v%�E�G�opR�#=�K�A�E'i��,!���{����G�+��0YA�s���d�t?0Y�cn�n���O�\�H��|���"e8w���}z`�1���}Fk�-���������h�(Y��J٘�	��s���u��_�����~�O�N;���e��b�WM	i����h�
�I1t"��q�R���gY�׾Y�Css����M�?�����)�>��e��Y����o���[���Q�2��[��܏�ņVNLF��{ Q��TJ����KW:+��j!��
ť,V`[T�{��N�eG#Dd�*��ko�!T]��c{N�`�N�Ä��Y�=%�A纳"�$�_y��Xb�BB�r��