XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����1�	Y>�9�t�3���������(��9y��gU��1�n,GO�7S9��?Ȓ�(�tS_����ŋ�'~�� C���^#k
����e2,_��^���-�nvy;��o��8�D����O��.����X���~�j��.�b�?�� 0a�C������σ�p�/L������y�}��%)�ʨ��>5�����$��}�x��'�
�W ��0�>�����Rn��ϚX#��e�	�#�zM��ri�`�OH��V�سk4�_���[>5�L�`�r��_�,T|If���!4�P8ޠ��8����ï�����Jx��#�T�	�T�u������_��u4P�D7_����n���7�P��ڏ���2d���k��LY�����V�=�ہ�@�V��o��#��DP��v��s��~>(���#�M�$��ix��oT��U?K�����wnM���#����
4lM'7�-����
D�L%�r��c��@����/ߣU��|����B�;d�G�O��|L��㖻̱���&�܍����$z�qv������.��]�aR�d�T����Y���a��PS�a_u4/����2��!Й1�/ݪ��>f��@">�Mӹ9�M�H��_�GC����ǰ$�׬W��Efa}q�*x��!������4BsE?�M�4r��=��4��ٶ�5vS0���u�і��j8���F�^BF�Fz-�W0ִx��D"�YO�q!�sm��حXlxVHYEB    1901     450��wN/�)<�̨Ѧ=�W\5�!�ܕ
��C�rY���׹s7+�s�V�����r��F�/65ۉ&��ov���s%a�a�~��>�4tP)k3� V��]�Z3���@(���}f��R�4�)Y�G�
�Ag�צ�`�>�>���$MȌ�c�t��� �����Wt�u֊�f�,�����v��pU��[:;�j�Og�,�7y �����~�j֚x�8��
��m��3�ڜ�F+@z�W�В8�%-�x�^l��x_��8LқUH�����Zc��<������'�>��;P���h�E����9Nƿ��\0A��(bdc�3Åց�x�
/�n����F�-[t���
�`�Ƕ�����ݱ���H��9$�t��H^��t��M.��A�a%LKSs���4>ҺxB�:uᑧ���9��p���{7{u��N�������7�B<���[����h��k";�'F?�-]#fx�J�6�5�ὲˎ��RKS�3x3�t0*Yw�֓���\����j �3��|�x����]�ѻ_}U�.��NWr(��",���>��3bJ0���[���\�w/UJu,��n2�+d;����8�0�@j�uX=|��1�\(�k9�z�0�ou~<���7��G��`��������O��Y&�?�^p�Q�Uw_�|5�)!��D׍N���7�����`�l����%�"�Y�ޞu�f?�+�?g�+N�0�q't�%�"i��b���B��Dۿ���%�#����9��^�6ț�ᘂ�i�qR�A�q\�(c�Ⱥ@SiH��K�㡒�'�c�Zr�æ[KL�TB�r�2�˚fud�]���PG��qљ�%��qc�mY(HV���m�B���ӝ�rG����(��'F�'.{����[.�o@�W6dL��G�up7:>�r��N��R����΢/��I>�[�Zৌ=�o��a�g9>������3�]���l��ⲹ�Wq�h�Ubg+C+��E�k��$Hru0��gFa�S�ޅZV��z� z�9���o3��7檧3��.+��A|�����IQ�a�,�sh���D
Z���'�o�����R ���y�