XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0j�{}o��Bc�6��~'*C�EC���V��d�|3�Bc^����(3����9P��df'��TA�����F(zv]���V���O{5���QB-x�ޱ��w
l�V6FzOߡ���ST&v��gy1��9���F7�;*�'K��s�M<j���q����8WJ"��Y������('�k�ѥ�(~?B��w�}Sp���m�u�j_#�In��M��xV�d��;�+i^ (a N͒P̄��y9�u���0bb_�x̯(ܡ�g �˚ �cDw@���h��C���7֭XQP����O-]�o�[r�����(��#�}*�>y��Y'd\���E�x�ī�L��q�<��!M	�ι�.Ʉf�g��u'K�3*��2u�Çz�}	�]��qѸ��Q�K�/���ā0k�܉���Sa�|,`�n�o)��~rLD�[Tю�)����|����e�uU�[3����-�����!V��y�(Vxƻ�g�(������f������i\M�4&�0QJ&��a��u������5��P�=�P�Yޘ({���ڡ7@0B��"s��5
y�Y��/O��D��|����[6g8�	�������� �q;�������Ϡ~�C���:����C���/�q�:7�)�cl�x+�7/�w/̭1��źV�
�s�[���Z��|��� RQ���ٝ��Y�$�'�Nٍ���ZC`��>ʯ�X�����G������8o�g�DB��wa��XlxVHYEB     99f     360bG�T�y�oSo�wre���I� vl�V���u�!��T�cά�@�� ���,��+�y)hj'�[1��캰TR�r��6p��&�t:��t�߆mwTŘ,����8" *�h�����DH��F��~�#�F�fN��E����O@H��̢���͋|�l�O�q]��1����[�������/J.!|���s_�,��av�;��6]��J׌S<�ힰ*�gD�ѫԝ����%��۠�m��H�V~`9yw`M�`���>>�Ć��Y�01��i�������c��:�7;0c*n��j�O����t�#�!M{9j���h�����>� �l���
0Ǻv�+G�b���G�|C"�x�����/}G��>��7i�d���B�mK�<ʫ�Y����w�N�&��γ�C�z�����S�i��H�\�3�z�Ϭ��8��?J'x\%�7U@>�T��_��:m�Z�g���&Ē*�}���u��#������wGae���U�O[.F%x�Z�
/��9��w�_�
��1�@_U�l�u��X������,U\�C:���eO���ݕv���9�9{��NlQ؞��i_Ξt0N�y��m��6�I� ������3Y�`3��*�0&�ApLo?�R	M���P�B.i�C��T�ŝ!�)�k�H�v�]�7g���n�8��<v��Wx4I�x�8���b7+ �A��%~�'��`oƤ�nd���Ck����� נ����Bbxs��E�	A���s�h��|C��݌���1�[|n�GO;����C0_��^$}!bJ�,��!���.\�@��_ Xu��