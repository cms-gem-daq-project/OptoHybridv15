XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��KB�ƁW�����6����q���|��\�r,<&�>�9�{���y���{�~k��\�~]:�Pq�}}>�]0��Ue���@����~�.�K�&�r��]�"�P�0K���kR����Q�~�z��O�[������0���Z8`5��V�abu�9߶����
��$J̶�����ů����dϯHS�����ý��t���,�j}���Lj��ϡ�	r[6��!s���g�Ƈ�j�b��:��B3�U���Dϳ�mA�4���:��1�m[S�T��٧5�C��[�U:y����t���:=��Q:�}�9H�(�`�=Z��������V�~�d�}r����̞�Ǆ~���O�3�mdSV��DY"xs9�g�@�zOp�C�������车��M9���|Δ��3eއ����.	�e����S�[�����X۷����x+I�i[o��C�۠d�Wr��g�!���O�����`5{��+7|��r?����o�6DU���JkD�sA_�(���G�8����b�n���	�YI.��+3ޜ�(��u��Jތ?�����SH��]�^�9�c���᳇W��������o��
��1�1�����Ą9��k���]@5�R|�Q�5g=��Bg
f�c�b��񏙏1�SR�5��q�D�E�YǠc�D(s�d��e��t�v�%B9#��h���݌y@�Ӣ�T����|�h)�c��u]fըW������GP,��S.�7@sXlxVHYEB    1d52     7b0�n�f�&B��!eZ�~Q4���̼���Q�%+���u�θ񭻴�w�%hpZ9��B�w��]� ��jK���S��
bW%��%��>I�Wn��-J  �z]jM]ܤض���Fq��1W��JT�Wr�p[eX�pLq����<,PL�aB�Ǯ�&n��I-�r�Q�����kY��%(z*֘�*a�$���$,��)( )^ppNi�֥�(g�8��z����̙j6d�r���s$~���{��5���hBuGS���zLs�쑥~[���^���F��ӧ4=�1�P1?0������"�
�5'^^x�"�'C=*�P\���u-��m���ڀ�m�R�K'� �YvA��Ó�������b�ƨ��KPdسKp_Q#I�u.��F^�K#.M�����1z8i�ad�U�	6�ٵ>�A"�"��|e��R77���O���i%9�&;$���?�yjL(pxu�eFٓ2b3����{ӭ�f���.���}z�-"�E�B�_2��7�������>�0J�lm�[,)3�~~���^��C[r���I>�|��GgK�n�
ya��s��)ZD��"�lXȯb��F�hGމ��;���E��bB��'���;�u�u�T׺��9���Z:H�q:5d꩜��qW�q��o�}a$q�A�]������F��N�W;�.`p�n�2��x;��!;9~j�����$��4���u6%��h���-�t�����7��V�&pP���sr@R*ᆶ��?��g�����W��*�a��vq[t��3C�w��"�Mà���n������/��]Te�ˤ(M�%�#�7Y��e�� �%P�@{ں�����&(.�P!2�s�%���}9��߽G�>�Þ*fФqb=X��U�1X���i��#%h}nGe��5U��O�B�k롄�BGl9,qS���M~�5����ai���qQ�#����E5� :�ȱBa��K��I�q�2sf�� \��� �6V��FX[�}�	�|��-#Eۂmʕ���J��澙��N����(G��p1+a23��W�8��u���jS����7!D�43Z9��j�z�U)c���
(3	�WIJ�|c ��W1�/��=kv �����J�ά���G$���"Al0�a�O^��Cf T�~CT
O'�+K*+�a���� ;���u�*�^[�
��U��a\���$�Eo����#�u=�m��l���d�����D�R����rw� ��z��R�]fS�nu����z���#13U��j�-�G��J��҂��e���EҸ�,�������e򡮪�:��� \q���1�M���ÇI&�.E�Ǽ�J���e��O��(��.�r�y�գY���o���ZTݞ�u�����H�R�ަ�L���pE�!Tݨ-��8y���c �zo�#@�.�ʤa�t�8�U�b�|�C�]A9��	W_�8�Y�n��� ��%��xǵ�Qj|-dقL+�=�������ӌKb!�j���x����B�~�"{Sp���|����9�Z�^�;�";�ވJE����7tHC}�ӛ�E�hDF4�=�a,?j�`c����^��Z貤B�Q���'ō���ڈ�Z����L��شA'o�pP	=�o��a6`Q��q�u�������ʘGП�k1L�����!+c�E�2�t�a>���w�K�i�v���Z���+5��K[�>ޮ�U1��ڥx��⎟H
��]���Ve��Y���i�x���>	����	3cc/S8te�����a�􊹄�G�>� �i3<@��{����.��0w6{`�^쿂�:�LZ�̐�$�(O�,��=�<��F�@@�7w�̴���Ӓ�H�:���)��|�Eq��G���o�����	��Kn.2�!Ն��ͼ�$���q�կ&�}w;�b҅�Qr���� "��BO��1��4(F!�:�K�!������[