XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��׀���[�ozdYX1�(5��*�9d%�:w�2���7�������GB��ȉ���<��f~q��ō��s����U�p��I_�����b:~ �];�h~y_��x��wK������'�"s��x߁<�$%EȢ6̟v+���/�H���c���M���x0Bd��J3ͳ%��-זDwT~����&��6#�0���@����Ӝ����e�`����[�
G,X�u@���e
��̽8���^�+?���
��߉�m��넅����&#���^֤&�M���M)Pu���N�5�n�*�v�V2je�{[8H���WPAI.�O�W)u�����Ɇ\��g�j���a�kw��}�����TF(��v��n��ub����s懶7l��z&��
$f���	�<Ҭ� �q|�L��2���b�w��,��!�>!a�I����X�>����I%�"xm���8rF=���sާg��Pukf���᪦(|���u� �txS�}��#�S�z�1zד��}�Y!���hcK�3���{�pW�p�����)�&W�T��p���^�fI@Y�|�y[&�y�E�K$*�L>T`�䛕��ǲ?�p"��O�(�n �=i�ը�AM�0R�������9�P�8g��
�a��81��o��k�B#%!�3����f���&��W�$TŒI���X%S��^|��9(�H�����׫���~���l>
�HjoXlxVHYEB    fa00    19d0sjO�jr!�(��)����T^-1L,���&��m��N�������,�^�a�Mܻ�A]��Ɛ��C�s3c}ȵ+��p>;�����J�Q�a����r���Iޓ)���c�:�B��=$;sU�=*�Ն���;/�ƅ�PI�㉭�k}�����#���^�:��p`���B�yet/V�=�mN�H`7�f���f��T��od*���o:��N��K�4�:�T���|��-g�A\W^Gz
��ұ&��m?�^�U	c�~g�y�D� ��E!7�aL���}u�I�QBv<��Zer�z|o
����;�TF�- ���R��v�S40~� »nt?U�����\B����.�ͣDN�G�d�������f��Fk�@ɋ$���_e�3i7K�}�h!�A"��R��]Q�e�b��v�Hӌ�q�]^�q���ճ��d@1{����5��E·" ��,�!�S 2����_~�L;��p9Õ�O�M�8���Þr�,<�s��C����l{�/z��|���U���C>Ez�̫k}����,�Ͽˀ�oUCzVV>{br�<�*/�� Zwפ**��c:��ŨvՎ���_��7���.A�q�$Q�ȗ@�a�����_-���̄���jB��'�5�4X����M�����鉅��,n�@�K2�� #�9��Y�"s��G�I8Wm(U6P}4�D��k�'(coa@����?��2O�K>b ~9�O��l�ɘ���[*����(��w�BN0LJ�����q��� 24��A���(�פzD�UZ�'A���v�G�Bgk��7���p��O�掤���*Q^A�D����}�z���K4ט�SEm��ۤi���tY+`�j�l5�Zf}�C�U���[e�MT9��7�����F?a�p�OR���k�^��������cm�K��6���R��Ib�!�|�<�7�I!�!�f�,o�����N?� �8]9�Z	��6Z =8���咰�2��hD��$�=�E�9�ixF�H�Y��T�U�w���������ܝ#�i�V�i�̯K�]�]Go~���F��X� �d�����)c�[�E@!�ɂ�W]�A�5b����2�N���@�{�!:	�� ����5W&��/���H[`M(�E�$�z���ې�w�����A�v@�Q��ΚJ��.����=��I�m_#��Ӎz��T��Ny����|��t`���p����)a*+����v��ʬ�I2�,�)���v �Ra�MKg�zB\3w� -�>��ŷ���]��A����:6{`�|z�'���V�w_W͟�i���(_��ּ.W.Tz�v�9;����jp8���qАe�
�����Sk��A��QC�O�'^b_�/�Z+�k������d/��`�f��������8�pα���e��˦��_)�� ȍ·�4Z�=��R��ؖ���t�������i#RI��*-�a���q���j�&Y*~���\ɳ��7x�(�%36Fn=݊�$F��j���#�a�;�~.6��ќ2�ZI�wX���7E��F[��K�����:&p��E���;%,+�8�Y9��rs�~�x��":7��K�An�P<_xJ9��抝M^V\ �����Kmy�>��c���6Q�y��)�L�q��|�ۂ�h$����ʷ�OS�`i��T.#�=��3����c������S.^
0JbkW�3�D`A�������	�?���ܦ�#<��!i�o�\%���1o��s�?�ܦ�#�l�Uy0Sn��1���(/s	��!�:{Pa�{���]�]x�TJ����O-dw~FA��ƥgB����tͨnfA���uQ�pԬ,�Y�� E�)�_Z�Hd��s��3��K_w�O�����\�;.�� ZG!	�W��s����� 5f��fBx��t]�߬6G�s����)֕KղZ�$n��49���G�#�谔j�ހ�>ar1�?JB�
� lf@�Yl�8d$��P5�����.<���ߧp&H��O���0�$�k,��틍�>���F|��.�J̕.������@+Uxp~�Z�U��f�Z��m��� �α-3���a���M_�T�w�@�0�.=u��k{W�c��9���%�5���4����o\�묧;c!�n�u*I���C)z��"j�_�P~��x���{��0�p���s��0�&��'�M#
��D��aP�0�`4���:A�$-�s)h�S��z�"ȭ�W�OA{@��o���fc�v��ٛ�)��
|Ja��]8�4L�p��.�+��Qf��Z����_����~=�]*X��swI\6��&L[����d�O�OF�";B�� �x�Q�1j������᧙>��{��f�CG��$��T�&��4s)"OA� ����w�ߴ�WL!1F2�6�az]�q��cIamy�����Fl�ʊ�Mm��
��o S��o��ŜuP,���C�s�4Yjz�lDH렍#``t�E��v�>T��5S�=�ҖP���tEE��	'�
���U[�\���Dn��'��7F"d9�8a#�\K���ff "����;�+ �`�=@�o���mY�W!g��u���YWRX��;��j� B�a������d�@f�h��2[�g�-�(��r���9H�A�z��/Eo�Ĝ�3�k�s3�%�-��� �Gg�s�Ex�t1�@�3��$Mi+;����qkI�s�,���R|��s	��$��] ��4YݘS��J?�qq�[zdV交3�u��J�$��R�� �@���\���Ht<v���oh^��棔�7�&ؕ�E/A�Y���Z���3$Ke3k�Ӥ��������M^�@Bʿ�+�F���TN��u�+�]��,�U�<��2Nc�-Ј/�d{RCNe���nS�N�wb;s�ݠg�qs��O���a
� 6�V	��<��l�Qy�t��wb�}��B5��1�oܰ�ˈc��y:E&�����ʳ��s��A޵�A�Qʦ�_���7�u��R"����H jJ^,+A�}��%��?~Q���wW�J�b:J��Q3�-�#�/E�j�?Qt����ӂ��8d�>���i�ƶ�@�=�>�)��z���`�Ǳ���R9P�y�B{��O{���⑰�XM<���`��D鴽 vŀ!!�E��;�S�?@S�Vb�硖{׻�1����?�JA�?�-���\�&?�� ���E��o��=��`���q���+4c�<���m ���6c�}��8NA�0�(���J���9��J>�>ݵ$}*�p���ck�'_�Ԛ[�]�M_�"�׻C�������]-<�_�z���k\Y�ڑ0���y�@���V��-3��x��=�cQV���E�cϑ��m�wjo�O��d��6��P��W~S_�bs�����G��4a\�4qDG�@`\�)�K���1��I �4��-��2`UT��ɇZ�.�Ú�4�"�SÕqɾl�؀�5�"tM9N�ʘ��F��YQ�lfؔ�@20^���c��$���>�����sT�\��E����N��'����������
��/o
�?�ry|7�m)̢�3M��9
r'�R�^,�c��?�>>�x�Ņg�����=~e�kQvm���7-�a��W�6qh�t�tG32<I�a��*��F��3�~��V��\2$��N����u_t����tvD�FX	 �qT��^E��W�<=��K� 1���+Fo����ӻ�m�{{�Yk�5�!?��^����lk��Sm`@? ��SL��葼����eÍ�"t�r`�?Kk�b(W9m�zWkO6�Ȥ�CƲNY�`�y)�0� Қ��X��ۃG��'^�	��}�>'��]p��GW�g:�q�TR��Om,{<휳�u�=�riCZ߮2��ZR߫�?��(.�'���ML��`6�'��*���<�??o{hnͿ+��t�#.'�tH�x�&�O��e%�,a2xЋ��[[�{�Z})=t�/D�깇���]m���ӄ����;-�A����*��A3}!�r==�>�ٶkԸ��~*�O^2	���q�b�*���Ť�"s�<p��E8 ��.^т_w������B��,��x`>/�Šw�y�wL�U���}���pM´U*}i����܅H�Z���+Yj�4R�z �o��)L1@�_�И��$f�"�^�H6b�2�R!��^�$��]hY��%�Y|7�պU��og�������Įъ�����"B��!�8���/�Q�׽ֹj)7�`�i��GΟS�nԎǮ��`jrr�WX\����g�,��/N�mK�"����^ʩ����"�d�W������Z���O�L O"q�e&V��ߕ�yd�	l�%���0�>���Um��5�׉)e/�L����G`_1�ES_{����ӴK
���: �9�r�%�L[yJ�;�����|v�&�#*�8�>	�������˻~�^]��w�c6���f`�G����f�?����ׄ�s_����1���t��_Ff_�<�%.�M���z˵M	͇#��Eq�M�L�m
z��6-$5�)�V��?qY�&,�z]��U��I�ˈ�����$��?n�_�&<uWk�(.]�����4��˩�_T��Mlw����?��#����z��&��h���m�"���o�)g�����
w�8י�AY}��0'Qpq�,�z�8�G����Z�r�F~�G���B�s<��~Cy��<���(O�.��q 9�Nu��B<�w��[N�����:�~2$��H4�m)_��,>�^;k=�z��|Rt��0�+��ݳ�a68�&�I��x�H�ܽ�/��l��p�4���q�^�U�v�Ղ���[��Y�b+��{�&8��(��� x�%-�4�/QU*��w�����q�2��o�1�]��A�ƻ��&���Ʋ�_1wn�^�Q	�f7�\�-�h�P��U������y@d��]�w.���rK����j)$�`9��:>j @(y7	X��c� �BL�"�S>���gKFd^������н�&r����1�a�8c��-��{��C�bز<�0�6�}^��y�T�毙����z��4�0�X^ەs�득,�|�{�89I�P�t�đ����&�	j����}�[g��<��V�l�YA�4[xrX�w��	@�%z�C�:׳A�����K#Z%�,u:b}�2�@l�j��?��vh��{��K8���-������3�0�C�c�K���P*���h�o�q�+9��b�kY�|tE�@���{^����|��;���ۅ�HMI������x���;��sΛ�A2Q'}�QW���}�r���]I,l;������.��_7����/�V��Ү�E�1W�]�;0R��#F�	������q�k�;^���6�4m��:���rJ�[��s�eB��?i}�@�RK���Om,�h$��
LȞ�ƴ�T��>�Q��#�)m����afe��=�\V����;��̪/�_L)+�tɇ;�u2p�(�뎈aPh�����_��%9�0�K�!h����/����f oM��kp%�t4����~Y�[�M5�
�Y��/�i�e@ظ�RZ��w�������-X�S㑪43B��{W���<[�.AJ'��;�g����X2d��[8��LA���[��\�;4��w�Ѵ�����A��BWH���lR,���M���H7t^^�6�5�Nb��GL9�aU�B�HfT7��@�cP���C�U�̴�ʃp"
�A�Q����O�G��
��5���������0��ާ(���8��7���=�a�r�j�1_��4�e�qs�dx�Mlc7]�)����v�Su ^i/}����Emf�N��U�S�OA(0��a�hB���ʼ��fT�kU���O�٥�Ǌ�TANö�y��� �2��X`h��dR�xD��QXP�-`5�~��͍N�&|��2V8�}	&b�nMp�3�Hs�`�f�&Ą8��:�^��{���|K�G �Mp�^�lęR�e����Q�K�%�K���4jHp�����Э��3����t���Q��P��-e���A�lv<�+�(k�����׺���̇m�@k��◧�D%�3a5���%����M7��P8�Ť��,U�N���`��>V'"MM�l������eh肢3K
7�P��X�D�)���d��[ĹX�SFpfKeM�g���$��潜��݊�z�a�P��.̡�LwmZ�g��u��жı�&Z+�f9��Wa+4�Y����ș	�lE��t^���MV���g� 沊-ĳr��=���`�{�3^&��3���w���Iޫ��J/L�eѡD�l���AԸ�U	̂.�wіI3�wo������WC��r���梮L$���hil#��2m�M�8ik7��C�Iړql�׾Wx@9\`����oq��mPj$�@���I0'�%�y=�tY�i�=W��p:�A�"�N�7�vXlxVHYEB    fa00    1630S�7�*��q��{�<U�in���l6��雃�s��A �&���C��B���6�qZ+��[��@�S`k6㫀�M#
��h�W[�)ԟP�ݦT�R3\L'�wp��"� �I�������l��������y����΍�l$��v�h;!��Oޥd�s*�-�ݨ��%�䴞kڜ�K0�^��d&�9�X��ґִ��krXR���<(_sm�bs�#|����ySnN��i�L�;с)����o�#�V�L�d��=�o��o�UքXi��*�Y�jxZtB)^��F�b�B0h��EÅ�$5QbcN��j�Mr oHM�Q�x�����	j98�����]��x����?���ɐ� 
A�0��Hՠ��������7�:��?�:1xU(II�p�n�Wa��������ضa�־,�ฅ��O?v6���D����I��0Pf����}���97ϬlOn$Oy���5̙��Ԛ0Y���%�Uq�N�=����_7�2m�#M�ZNJ��|z��l����-lP��V��	
�B	n`8ßށ�Qٗ�&wϼ�4*������
F��ퟮ�C�bK���u��p%�hT�*��:g�[�&]L���J�Ɨ;-B�j<g��g(�ȎR6���a����N�J�ʐI��+�����0���4~����:���5�� ��iJE��#zX�l3�����cu�X��s���+Cl=d�ǟq�@uX<|L?d�Vf�6�ܮ^?q�@�Y�'O�ܘ�a�B?�Mէ�z`�,z��_{=����`��/��7��ݗSF�T����`��}]�f����_M�����9��W,�-{�؋�gŔ#Y���s:�5]yn�<�
��:S��<�o��uU'u�̭T�Y�򰋞���靳�H
���6�C��o1n��
ȩ����[`PUZv�5��]ɧ@��U�r],��{��]�Գ"�'	2��Aň�����\`��2���P8�u|��,�w�y󖍉3T�;<�@�u��x
z4��!���c�
n�b�MaA��E[�C�P���s�PZ\��� n�^�Ʀ�{X����8���C"��T�ȹ\���V�����#�2���INͳ[�T=T@i�W��$��e�z��E*��)��=�F9�P|l&�v����<���_�\�0���&��̨��f~�:��b�X{��70C�?���0��CJ�e�������w��hf���_���J`�L���)�:��1�,�\�+o]�L�/����B�⢞P�;�Y	@u��8�ԚNc�K��\#�bF#LpP�G+�7�Of��<3��7��X����qƃ+���|��W�e7���Q� S��E��e.��hi���HҠ��霝 &���P��rw 
U��P
5o�J.m�LN����dʩ�b��|A2^P��ei�r�����J͉Z�9��wO����m˼��؞��|ÿF�Jeq���K>a�A�W��Kc���0E.Og�{�R����H��p���Qi{�f�޾p2Fz[�Ҁ��趫�<�����B�*�,�{��N�6���W�GYAp"�KK��	t!� ��'�=�N�p@����p���@����l�����N���`G�
�6Q���Jhx�0��b�r���@��e��ⵤ#�G`��7U,3�B��;���=2z�N����иH�)4SO�nT�X�x�����7)i�#�f�S���v�GOi���rÃ;�%`�[xoZ>��h,Jr萎��V��3ޭޔ�U�#��P�­��\�c_�(�04�e��C���!���9�.�D7�E.����e���wx`y�km *�S����t��~Pr��V�L��d�#� ��O�+si�r��=o#(����C�^�^q�\65�N�F�c�īN��k�b�������o�2��������3wߢ~Z�S]��y
ڊGd)�K5:�eN�ļ�BL���������$p�}�]�"S�֨h���K��#%L�Gd�x��&)��� B/u4���c�Ɛa5L �$��g�K��=A�OD3�b�
�7��VQgt�R���_�����:,����=B��5�%	qψ�����\��K�D�h�^`�^���~m�%��	��x��*�H�#̈@j�#�<m�$�?��@b��w���Wґ�Nf�b*��?�����w�u�+H���FuH�5�y��H�lK[%M6������W��PN=�ư��p����Yy0J���ì!GI�i���<�O���+=�'�(t��0FPb|Z��Ｊ���X���H ��?EY��	E��K��b�U:�+��:������J�A~hl��ev��)�N��m�*ƍ�o��T'aDV��/>�1th�{�RJ��޵$Ң�54����0�X���1SJ��D^�����c`&�[g��� 7ϡ���mx\/�m{��"}���W{�g���Y&K*n�x�w('���1�7�+hۓ�F#D�f�B6�j�T�P�˦d���C�&*Pˀ�-�ndEl��[�'��2}L�_�]c.$6��U?��������,�&i���?g����Y����F-p���|uB\(�'ϩs
`�C16�y�!���m�*�S@O:N�\�����M0��I��|d���~K����Hr�|����q�u�k/E�W�*tc��h�2�jE#���ݙ-F	]��A'_�^�<ޖr��x�R��6AR��_�wH.O�����TƭZk�閵�2��L��!s�:Ĩg�@{o0�ZrT�o@���`5߂��l�VLɏ�-6�y$D[t�7�����x�)"#�-+���Vz�C������& �,�@������:�|����N���L���ϡ��3P��Iy��~�w,Q<���;�S�v/AX�mi��?���ZB�*��u"'��ϑ�'����IK��<��^z�S@�	׊5
1w��~-���CR?g�wa)k aK��5�����j��V�}az>D2)Օ�ῦ8;�U���,�K��U<�m�4�f6��Z��X_.u�;;�+����Y1<�CEq���4s��W�fǚ����"���l��Q�>��G���G����S]2+u�1,XY3����?C0����I��l���*�CK��e�h��L�0�%`��R��F>"�]�'��I']`���;��jC]�a6��'ԡ�N���9̉����{/w�q��H���x�>�㘓����$�s��4Mo�\�G�H�����>�%ә0��z�̨2Q�P�O|V�E$.B�����B	�A�8�s�|��T{������^��9�	s���.���M�����-�(�K�S�Q(M�o9�>��׿��*�q���P����Vܫ����թۺ���{A$��^]]����$c�8�H���5���*J�e&�>������/�Gh�һ�u�s���1H��&��`CJ�>�3	b���z[؞�VT�:�IL�z�ܽ�';����I�Lo�*#K%�p�|�G�?�1R��a˙���4#�'p\1��2��w� aYմ�1�B5�i�^�C��z�˿}��6�n?����F<#$�	��������wD��	X�
tD�K�1(k��z����D�-���\u��(�m7;�,���s|�t#voK�t�]��-�B]��!TO��e�O8.��B	dM*��r�s9O�_]^2�y��d�KY���~5��Ϙ��i�s겻���'!&��6v��Qf���w&�۟�uo�B��-;������Zj2eiw�.���
���$ZQĠ\�1<�1�:&(�k�H�`o���TB���HyIj0�Q�v��Ɔ��i�6����M�$����랡�n-Dl��q�+P��K��a�P�ɍ���W������ "���]��M��Z3�0�d�������+�[(t>.^^xW�Ś�@pG��#-kp�:��;�4a$����x��B��ѱ�z�
��2-$�_i_�t�����F���WUaTL�W`�'�S�G�c��1cН8M�R�&�{�����C�21pe�i������V�mlzg�1H#��̌=����1��2m;�kE;�y;>̑aDM��{���J�b0b[0���k����#���������x�^Ād�V&�'�AԼ�����E��ߜ�Jt �$=���a��
9#�D�)(�|ލ�������J�Qi���z��И'�	�V�/�u�3$������;D`�ir'�ʞE��ϣOB[P�m�� ���/1 گ	QT⃷���\d��G�Rl!�+.c�A��ǂ�vVs��t�G }'Gnة+8�32(�$j��>���[�Jm��}�U=��\��b-�m���ņg��:8��(l���O��� ޹aËW\F'�o&�V�W�)_�g5(j�v��;�2�'@�(ݢ'�� � 	`�A���ufy��Z�ŵ��:��)Xm�[��@/u�����d��N	Kɏ;|0EZ+��h��2)�!qXn�!��A%�=�$zh�`�V,�sM�A����x����QϾ?��Y�t��ER�*�%�'?�ݘ 0��o�ϡ-�7�31��{�眀��5�T��6���U��]�:[�I��a�ҔwÀ���� �i�v�p�x�`k,:�n)��)<��5+_�6ݏ'�f?����至J�k��7Bf�,ys]��Jz��h:��WeW��)�E�M���m-LX�o��*Α��ۤ��6�2/�A��x�L�a����k ��LM���_Y��\�yU}��0��<U~���:��?;*{�*1�,@��|Ҕ mQ������2W���IzFM𮺇ZH����2�aEr\��(��(�#ȣŻ}��|0d�0�Y��C�<���'��(��g=��*�i�jk�fD8o����\#�^t����4��UwRg�jN5ԴS�B����d�|	��	��!0�wq[���jʀ�@F�n·h�����I��䠰)��"�������s��Ȭ��RN^`<�0L�ٸ_��m������_)�x�ͫr���[1���u���".\|$k��#VZ�U�)������ϛ���6��|U<���B�M���J�L�Y'WDձ>��f���O��;�� �-�?@����J�3M[Z�F���?cW�oL�>��FR���dY�}��on����Ә�y���rQ��R��NYZ�_�c���X>��)��9'u�h��S��נ�+�x͂\ s
\r7�.��&K+	�r$��=�$����4�@(�ZGs��� fz���l�$�q��<T/��UV�'Mv���B(����("�^��b,&����衪D�g�h��ۭ�k�X�3������t	>�22�6���)���
qk���p�� ���S�����v�6T�uq���Q�:J�o�#A.�N�~���������ڽϑ4�OޠG!9�b����"��[�\��Ն�j;$	E��i���|):��V{ƺ6�l ��0]ͱ"���qD��LOy����Y�K59�z�I���)�ҹ(�O�r�l�HG��Uk�+(jQLݠ-6�0�V����+6�w��u0i#?!��.|��)�����]�u(����M�8��p��o�%���뀷���u��YXlxVHYEB    fa00    16a0If����y���x A���?�|�'&��D�&���$"�t&���XǃDt��ˣ�:p50D���}��T�P�6Κ0��},���]��4�yb�d�=�{]�X3�`� ;���vmj�{pk����õ��Zpvo�u�W|��&��F�=^��Պ�^���<�3�����e*J�e�>"�7�32N�	��H8�׬p�����<��t9�ȱFm���� ۿ��1*���5��ϙE�IA9�z�}�9}q���s}��?g����m���@�4_ŉ���)�A]ǳ�cO��^�΢���IpMev�1��6v���~m��2�ս����%)�'&F �A
lϸZ�!@f���t�5���夬V|Aw��L�.��o�EI{rc�K�/a	9�[JRɛ�����3�۔��.��3�4�fy��`�6�`�Bs����W7M��[I�o�Q�����+�($�6��ck|��WmZA��g��<�"��RxR�"���y=<`�~�kӭ:8�m?�
��������<��2@]���EJ펋Km���e�'��f��<����;3[3�n�N�m��ư��%�M���~��'�����|�۸��T�[�������U&��Ӧ ^��T���XԜڈ��G��S#��"˛�.����]o��Go���@"~��+�y�,���/5lC�>>ل��.C�B�aV1��bK.�7��.ך�(<�C2	��i��,������:9_�\/\toh�7n�MD߉$z�z�U�~�'C)�A���u��楧NeQK Ƀ�6��z:���?�H4������j�*t�������^�v�@�d]]؏sԟ2��Z��t�oj��lX��TO�r�`��:��)M9���$���/�(��vP,rXZ�K�aٯ���MeW07S��3'�Jx�!����k�ݷ��ȐJ�~r�v4�b�}��<S�tt��=�����Ml腤	�2a� �IruS_��T�����ߕ��>f]���s6�ۆ�K�:��g��������2�FkB,�6{��lĀ���nt#�j�Gy oZ*E���z 旺�c4�ۈBΧ�J'~��c.�q�CuP̧̛2\����_R���an�l��t�#�m��8���l�*O�?0�U�z�&��ƀ6@�y�e��BU�][H�����k��R�����Z��#�y��sy��V�A!5��f�@�߷rw\-ck�ѱ5fY��1^#��T��u�eź������9n��Bd��JW+��W��ihp�Lr�m�\��3�c?�
�~�[x�`�(�����Ao'��h2��v�������dJ;4*
��P�օ��y;�_�>{Z��T]S^]Y��\�0R���x����^�W��Z�Gz\�u@�#�d������/�z��w�!�d��N�냎�j�
t᏿� }A�
B��Ց�ALg�x]^��� ]�F0eQ�+�rv��]���@cfA�����&�yiP��I�E��צ#���a���S1��R�����ApU#��gJ0�x�}k+�*��*U�����r�$[�0\�� �>I1W�'K=K�n���i�+�I�����j��J BQg��j��q�����-��ԧ��[���.�&��h��LWboU�:���zd�4#�C_�u���m��:ƜQ�b�m�Q��e���e����?=@���S���h�ő58a���(��C�'���d��X�n�b����d�A�U���.��W	E^Twϴ�j�TPA���E�Rnͽ��|�"����v�����ͱ�f$52�=UtΓh�1���&�3��K��3��}]`v8�t��y<-�[���lH�e���/0R�c��S=@�D�43��.�4�<mn_�/ӧ47���M��,*����b&I�=�4X[��*r:��ک�� ]mr[M��䉒����j=.�w�nC��6�v���Ys��=��q�wOlAz�`|y^0��P�w�x���Se�E�������>M$W�r]�ҙ��,'T��}�EY��i��P�n�ou��ꄴک�^29�	I>����<%,B��LTB��&B��8���{�}-1	��݁q6����ďj���faQ��j�P])��+z�<�ޙwV$Twm�f�w��7O�lW�I�$���9?��Y��uߊ�:��^�c	����X�Dc-Oj|�A7��LTY��n����M�\�m���r�Z2��TT3�����(?����;u��f,����~�1��P}<y5�A�oU�����X;��d�1ne�K^���$�e]�����E��^�k6��EE��M �bT�W���Ϋ|Y?�⃥=V��/mB���Π�t�ӵ$��u��ews�ۓ�����-aqs�]�������I~���,� �z����>I�]V����O���6�D?3�Я�S1WA%s�M�xw3⿝QŔ���H����<R墏V"O�*Of�8�|�moG�(2�C��[���׏�~[�Bc��#=�Dp/��I���(��uƅ!�PyUH�����3��!��=�{ �-��!�М۝�p�6�&��T<�lҭ�/�H5Ї��K}�FecĲ��g��4�Wk����5���0��Gd8�|}��<k�[���#3�f��烱���q��#�����I�5���grX��#��D��H MC�`��⨴�c�)~�Ryӭ"�EL9TL�k�������)��W�7��^�7��Vw��b\���N�?6H�!�^?�v���fሃs֞�v�K���kF�ąn+'x&K圜�l�<��VHv��A��׃]L�gh$�5H���\���9���p�.�Kޚxa[�J3%�p��C��e�
/��@f��6k���*K��������^���9�B��#z.��Õ/>j�q�T4�skc˸e3c.XL0��V��M�y�=�j�P|�ꄜR�+�ת� 5��*���k޴��,wwQ����N����DAu
M�\pJ��	l�F h/�RN\cy?tݳ�_%a׹���I��M+��V%��@�΅ۂo[�Z��yJv��d��#l����@�6�f�E~�~;�jJ�Bħmɇ]�Sj���L:��^�_?*BY2�9���|�G�fD��,��
�����-�m�,wm�#Tȑ���ԝ��D��鱮�1�,��	Yn��ۧ�U5���%gVD��T>���ࣟ)���U��G�W�I�Ty�=��A�P���6���)��ON݅{LƜ��!�5���r]F������͙
V�R��U
��۪�4X������'�>��s֗��+q�<��ev�--rh��?E*�xq5��Q�=H2�E �ӝ�Gu�8h	F��������v�����dÁ��A�,�>��*��, l�h0/M�]��I���bD�ے�/]�仺���M']J����5��">2u�#�f�>�$���P<Lg"Ӎaa�w� w���NN!��f3,���D����љ_]�����/�i4�+SIB�~�G誴\�3
����:�dԤ�r��9�P=�y�AS��f��� `V��W�<\���Jc��.k4|���b���0�LH}�u� �m�'ׇl���,�6ӳp�b-���Sߖ+h)�ʜ�l�4�_	�"���,͚��j�pЁ9���&�k����X��,�� ���C~a�-׺�9�3;�f¬��9��Ci�|���n�x�FF/U%��"�~�@�v\XsHq�O��`5'iL-r�F��%o���\Ĩ�\ba|�y8���&���8�G��|ނ�gb8J^jϪfѹ�"5�
��cr���=���SK`즮H�m>�wp�����|\�-�Bk�G���~�V'?w/�3�C/
%��
T5�Bi�����_��2���vG72{=�JqϢ��}��+��=�f"�v�grV�OO��0IN��*[l�~˭��M����l�ŰX7I���{n�a'���+�jG�Ԇ~r �~���8������xGm: VĨ�������wo5}��68�D�N�]��Յ�=��t ��
�_/�:�|�5dL��z+5�D s��� �'���O�'��t�dNm��E�(m&��aoN�ITO��3pB�]J�l��������VA�H���^��lŕZ�_�<�l��n�P�pZ�dΩ�t���)��=9���ސ7S��ԡ���,�T#є�ϸ<�J�?=U\��{;y��ZNEjH��~Ңt�b���.Փ�?�̈́�(!�n'�r X�h
MBi�^��;[���e�ؽ �]Dg�BV�Q�]�K�ȇ�Ө�k�\s���~%�0��<�C��|D�{CE��в⡈#�����s�
Err�Uٸ��ed,͛�G\�O��d�>��,E-�*s�sZ�*���lPB*e�މ��j�?dG^}�A�}�Q4��f,u����߻�a����$�����e� ����8��� �E�
�G1lF���g`�b;*k>�a��#؂�>�3�y{�e���&d�S��3�qu�1�4��r�B�cԔ��Q�s��Н����^:C�Gy���Y�	c%�@�¥�����p�iu���>m�q���p��IUT|���_�1d����~��0C8��OP�U��i!�IH]� �����!�*�nxIo��$��Ԓ��Ə��6����"�������=D��+{��W��k�5�����LEY�u����jQ�Mf�6ҿ�P,��L�?�C�����ZSu��d���`����@���rê�"g~zn��hrǍL���&��R՗���3�>Ǥ�Y�B�S�A~�� ��S- ��1B�����Ln��)%�,�^�6��L��YXI���ax�W�@+�������o��L*�zm��Q0���z�1f�C�j��#H���\mi��J;^���W��'/|�<2��4������X?����D�~n��q���{����vj@�:@����AG�Wb��KmW�mb�.N%IM�m'tCk�:C��	�HZ���o�@�T8���2Kk{hm
9��,`��W��{p�r����b$ݑ�|r?qU���m!z�胰Y"��Ҟ�U������Q�!ӛJ��o���%��h�P?��c�oq˘X��1�<����y��9$�A�V䂣��Rk�5[�xr_�@�Ja�n.�eQ�Eϛo����!�m���A�ڕ��*J݋Ie������r�}���i��b��o�lv����<m���NG%2��u��L�!e	��d<H[�"I���ܔK�܎.;�l;fڢ[��_(��ߧ�����$z���/M��QЭ�����3��+�����ht�v�2�}OW�2:����n���|ײ$dGUʂ�+��?O=I�׭	^g�)AL��tT� ��/ܵEJ�m�Ͳʉ��fcO���H��C�b��+|Gv�������)G���H�����]�UIjL��� `��3�%��\�CQ�J�7��A�q�_���|���)D��w����g��.�\l�D��tԴ����[ȇ��	@��flT��z���Y�����v�i/�Dw��#�6�q� �!����@�!�(56�6�i<���������yޏ�x����a iy�=Nz�pcm0XlxVHYEB    2889     400^0�݇�wi�%��)w���BD�o^�^��}*]�9���tD��
� P�����Э�4mF�ܡ�1P�8���<��ݶ �iP��[��*�z�iZT_��������}P��U+#T����\H����	�riQ��:	߀|L{E
��C:���.f���m�N �y5����Kv��Ԁx�a}�:����f���[Pb0�3�Y|#�	減��M	v��߭GSLޡ��[��0��P��8P�	�S��5b��A��_�6ߧ�^6������#��m�I���B�p*�t����
��E�}>` -$8�m�
��:����

L�=�S�`סm"k�	,t	J p���g�R�b�jߙ�o\x=�,�l��:�yvґ^"B��tJ�]֯��$W5X��*�g��Z) �'[�_��@p���Wp��~��q	;��[�{ɲ�I�u�%�������C99;=�"���U�#|�%aВ���32���V�b�
*�]�1�`����p£��w��}r1$�|���~^ʕg
n`�g�c�a[�W�����H��$#��/��{x%������ꦷ?���U��,���k�&2x��ƥ�R���:�%|�Y�#~���<۾h��&�����䇪 FEE��i�B<��6���͠A�����B�����!�-g���2�s��U���l2?#L/�!1��\ރZ-�>���VKfn<0N��Y��6�͍i3��i���?�G�]�]}��}��nɘ5e�]�8��f��qB��6zQhVç<�+������B����5zO����'�	�<#oǀ�z[�N4*���a�+�ʹb�P��U���(�h�g�Y}�M$��,��yټ`�ҏ]���/-���s�{ۜ}]k�j��QaŐrB7X>k9�Xm���E�;x��{�%�<��ۧ�U������KpWUu��u�����.ڿ9�J�*7+O�z�ۍ#�W��+�A�0~V;�2c���dl�tr	�+�"{V���=,Bf|