XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
D�s��h[�VA�"��"{��׀:�a������8��J�(����2b�d c ��*:��{��
��2fO*:s�
�LC�L���J�2�\�#m���]����(�Y�J�o5�+��:� ��vI��.����U�>�'����
�>�O�wh~�J9[��j�
qU_�����@S9�bL�J�
����䘼NAW�U?Ea�+0�F�G৘n��}y_�S��7�����(���\D��j�7b���*?��xK�� 5<�x��e?���)�r)�M�8?�fvF��\�f��c�@�Qe���5�8r<�Rq�"I�H���}j_�D~���,�P� ����q��[��!�{A�!X�Z˩���)�{����ǓWW��p+�~�d���OʲPjT5�e@�=X��dĐY�����]h2�� �I��D�o8���Ɲ���%śekU�+q��X1Q�fW�Ђ�����)����
�c>��'�@:��C�,� ��P{ܠ gjݰJ�N�� �ޱ5�D������!�o�-뫑�J�:2�H�v�w��I�̱�k#��~n�^�CT��%�'����f�[FG\$]s��#ϝ?o�a+-K��i/T Q}��.�B��ZY�K�޸���*�2Q�:����T@��O�����c���U�wI��z�Q�Q!՗w9��;����o��;?m�!��s�(#�=�1��q��c�[�a�M�{,@���P�J1/T�u{k�L[�sV�<
~�
XXlxVHYEB    2864     8d0��-H��C�;4$s�*H���_8��F��?�؝���ɤc��`��T��x$1K�x��3��Pa��_$��dS;�5�|pC�����G�#�g��Џ��.��I�ܽ`�YYKM�a@��g8����p�Hf�e�LA���ʷ� �uhI���&�!$�#rT�>ܿk���t9��
����b֗��*kIj�����x+g'�A?�bT5���_��=��m�s��MH^�� ��X=p��@���˿J��O�Z3\c���8ąKeM5�</!��U�63�ht��;�%ef�ZY ��S��9�L�'�h���[�t������hK{(ۦ�C��?�j}U*5n�B}�P�|:�!w+�=�0ܣ����JiU���2^����lLݍ}k�d��7��)E�#�*)��r���t��R�	t�D)"�T�u��j^���\u���J(�cn��~�Kշ��Β�-.�e��G�,b\*����U���l<�t��O��E<�sIW �21Gq�n��\Lk�kj�ZR��� �4*���q����LV�$q��oХ��
��%� �u��zWq?�_hߡ�	����l4w�C ���p��%m{��h�8:ҵ&�8�����h��u��G�<75P@�
��l�U��v_L3����-Q��5��$�l�/�Ohs|��W���	�#���'/��DWT��Ӝ�RjEgV�K����Z�U&6��C��]�٘J��9^U��CSXN�sx�M�+�ϸ��%��x�M�^��e��P/]�����B"E�y�t�p�ꊦ�	I�Pe���9��<n1�j���)� DZ�Ad���7ٌȟ���J =k�]���¦(�N�-ЃF�OH㸝k7ot�4<���t1CI�
� )8�$_D�����2��6-*���ON9�np�jY� e2r���w7��@���s�����Q���g��×̌{T�yoV�5R	�X,�:]�?�1��P�ļ��H��!�ե�*��A1T֎S?j�M/�k;5�5�9��{Yar�r��<��;��0�&.�T��d]�;�7-<AFl���g�!|�^�`��4Y�}M��r�j�K��f�� l������n��}H�m���B�J!�+Ɗ>c���t�؁�z�!�l��P��
�r^�:�<��\Q݊_�$���R�-��/+�3 ��K�N!���$QRIg#����M%Mu%�&|�}�Ǆ�ՁK��S�t=�E������TP��$P�}�J�J*�b��B���f�0���I��qKa:x�X����%��C��8�[D�vҐ���-�hّ�?ם��#_-35��lr.�.Y�,�W,�og�'�;��؟���	���
�q)0�P�I�����n7M���G
B�,�(�=�*� �2��yy��H?�Z�f���_J��gf2��Ou�'`$禼-;���^���r�r�] ��10�]�7���'�F%0��N����m��B�|��lHs���ÿ�V��d�q5��_�Ua��) j�?�Pڸ�201�f�v!�6��	*�`����}2 �3t�?�$�e̪�R��z/t\6�z(�v?1 /�,A�=���j�H�7��(Պ��w�^��I��	�	!`�4�b�}X��M���i�	���3]]���{o���ؖނ�����W{w�O�RT��\�U}h4X�͉x��;t@^ۏc�à�ԙ���������l��nAe���l�ߚɸ?V�1�ý4]�I�R*$�fke�{�3S�S��o�2��b$�ԋ]���n��:F�E�K��<8۞P@u#���Y�oޯ��������uMyܰ73%��l{�Fk���)C�àQ���w�u�Gi&���e�Z�E��"�������.*�Q>����n�]Y41��U�>[��ۿeWR�1o�C0GZJr�Z��%%��f���٣b�K�6��"u��W�V�b�+̖�
6����~�i���ᵐ,5�u^��I����5�5PoD�n��.�q۫TP��ب`aځ2X����;��򛆙q��م<�}�Wb���ɃW������g����/5�RMb�Ų�T�ʘ��Ի��{Ų5Q�qNd�hw�/5�m���_�6�+s��/4��GW�+�N���s:��y!�h��*�gSL����$9S��!xN���B~p���lF���~c슘��ҽa2��r���`ʝ.��j6"�E/Q��A����