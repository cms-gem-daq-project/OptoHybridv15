XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)(�b, \/H�O٦j�̈́��Q�;���
�WC:���^�1���^u��( ^��"�7$?2�siPIH�1&���f����W���i!�K)A�6�`�'p!��c8���{"��6�VK]���vz0����0�]R*�*��҅�}�hI��%�}t^p|�>�m.|NB+I_\q�V��6ٵ��]�L����������[�:5�;=i��O�;��g��.�8��7�߬��+��_�����6���5�5L)(��u��X�D���&(4�3ퟳZϦ���s�FJB&8@�?����s��z������*�� ��i#�I�a�	�����[��:R�|=ڄn�� �&�^X	 
@Z���גY��z>�������[1�W]�(��O�z^\CIDEZ�V��g�]J�7����Af*�M��0H��繬��s3�}�kҐ���3�ܽ���?|�ҢP�A���T��+�[�Yl- �>�����a��ڥ+��ao
A*T��>���e�Iy�\8j�yG#f|Z,s@�H ˒l�c�wHa aN������.>GTx�����6�J8/b��� ���D�d���SCˆ����"�;p9,F�����REpx$�Hb/vA���K�K�%L���*�;�`4?�ɼ����C?T��h����΂���)�m?𩙓9`=�W�{N�1U��̖����ףb2 �"�R9�!��I�.�#�8�@�q�p
]ғDޙ&
�<��ͣXlxVHYEB    156c     590�9�حr>�X�Eև������B}�WM�l~�yK��[V�1G��S����DO�]]��&֊�Aظ+���ɊĜ����w(��&��=�g�(�c��HV���}�.�$uaH0*I�1ݵ�����t\��M����?��@����ͼ3yg)�<�I.��	3c��T��덵=%��n�(k�q�|��Cɀ ��"U�`+^_��ggR�����H���ث����m�
��Z��;�B���(���ذ���,�'��A�6`m�7K=����!��(Gj�L��4��Ռ�&C��cN�g�,�:��܀�g���j?�o|ne oK�D���8���4��7�?�ݥ����B�ĩ��'�g�����C�<�`�k=��l�2&}i�#iN��1xM̞�E��0��ZWRzM�%p��l�j����ې��-�Į�d��+ߗ�������W�d�
I�!�Iu<7A���k,f�1);���.M�th
0����0�nE�*��Ae�_�"��A�'���*�5$��F*�6z;���N�m%�U��艙@�:����z������\�v]����)1��k�����'`NtSc=Oɺ6���-��TxW/� �"�5�Q��)�)��'e��N���t����޴m"��V��@3�/��S3����n%�R�ZP K���f�Cؚ80H�%�p�M�7���5Eo4~��U��n��A؇�� `��I���Cئ��7�V��jo���@n!� �t�L��1">�^Vǔ�'�==�-r>6j����kO�9�����+����]���`>y�``Du�v���gQ�s�biI����̼�E�F��=n��.2S�#z��9�������[,�ouIan���1��3����fVb�%�7п�aD+��������T=��H&�&5a�	m���S`�*���:��*�݊�ό�&8����� ��hUMP� |��}?L[^
�xs`���I@!&�6$��Û0�����ٷ����K�zHh�#�z<��=0�h��Kj|)�?��8!��t����檹�ĵ�R�W�I�d*�?�uT>�fg�^y�Aj��5���3�y����Ybz����A�)G��3�% ������Ͱ$]��C��Cvb9ꗰA#ƶw�\SK@Al���郕YXqLXY�e,�wP��&HL�H*�\2O�Rؐ�7\��B��Bi4��"��Ww򜩲�U�5F�]w3o �6��<R@|vNu��RL�p�r��]Pu���] }D�YM��l.�,3�����>��E}�p�"^S�Y֦�����3��G��N �0�5�֯@`V�-�եW��EC�|��]�H��%<E���s�����(�����I;���y�B�Ώ闒�3��[