XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-m�� u�:���RH��ʷ��{�B�b&�!?TU�*��~-C��*� ��{���@u#Wc�����X��/fߛ����J]79'�A\�1G�����%�Vπ��!�o3*vM~Z��I(̑Q�vkEa����N��ON�� ����wiXa�,H�ڛKe
�T��Me�[���û7��׾ŧT���!�ݤ΢HG�ea]�ЉET����5��%��Y��}�cΑ��;���̘"�J�+gx�ҪJІ����>��D����R�d#�'��I�w����ZƜv��xҔX���x^S]0�x��P��zcF�����>����b� $�Z��d�Zc�]M(���Z��B��u���(��ZZG�6�C$KF� �Ϝ&�ނ�-׭���\�J� w����x�f�u��u��7P�ӶS���:����]$�x���o�v�=����|�K�ۡ���ߩ�
V��K����hX�U=��^����|j!��y{��i1B[)Nyu�!b�ٶ;�=d�'�6&��q�j���a8����S�~"�5;�o����&��ܧg�%-U������9(K�xJJs:5��U���%�a�V��VT��=5=UQ�ì�kž��MB?��D)��i���:�� ���f��Q��%o�E��������ϯ��'�2~]���|0ҩ�?�w�h�Se�Zx&� j�|����s�٘H�n�}�u� �B�̛������)���Ӓ��H(o�����rK�4��p-����fXlxVHYEB    2695     680�1׺�QN�n���E:�X+.l���o���lS��r"�=\�'��&"Hz�~�M$x�'Q=Z`��1x�03�p��=�LL]Lړ\�b~��!o7j�G�m�h��$�;��Ln�'N����S2�(�t���rS{����Q�
�MNh���5_�h��\q�k2
���茁�4�[�ի�����U��A����.���%�>�V|\�&�S7\A�%L���6m��Ȗ�_�o�D�$x�}��4e���Ќ�������=�˃����Hb�;������.��S��@��ܚtF{y��85�٧|�*�����ܭ�&p���$�݃<	��[Zm���_���Ң���z��lԎĭW�`��6Ͱ��u�O����Ӂ�r��w[����=���U��RWJ,���,�f�e���oĀ�c`jQ��ngI�~��G~�r.q�����)��w��� ��u��S�}�Kms\a���"Z9�>x�����n��X9ؘ��|7�1���'��j��.-�5x���3��U}�vVؒz���(ot��V0���Ezȑ2�4bsh����˲U�-���Pj��*X�5q�G���㡤{'�"]�3�ٟ�E��T���@2�j\:,�݂�{�:l�i��u� ��B䱙_&�vK�J-�Dψ}�`"�"�%��`�(�}┄�'7�Ri������)���G��W8����X���h�!�[��M�6�POoS�4����}�^��)j.W#ш��9��O"��Z���0�ٻ?������|<m}�P�J}c6�m��.Ђ�����	ؠ�\bR��q���`t�y���r�t!ck����Gjvd��}<���뽂�!O��j��_ZI���t>C;o'�,A���F�0�=6ZAX*� ��Ӹ�V�ֹ�<φ�:���԰	b�S�����JB- <b�!K/A������r����#o�>��o�WPv�7,]�.�1�����1�:�n� ��d^$�Us`�����ϥ��k(����h&_k��4YQ8�/ds_n(���ӫ=Cb-��~���Cl�O9�p2��ED���+Y���=߸��$�?Ce3�h�<��(\���q��5��79֙�t�Dy�y^�``!*��q笎q��U���6o�9a�7�"�.E�ٟ~��h�\{$ƛc��׼��G9��\�9����.�ʩ)��u�T���F��PC��b��rӖg
Z~��ژ�F������X)a����Ei��V��7�ˠ��T�o�`۳~�n�{��`Z�D��>�	��D<~�q�C��!t�Pջbw�����	-ݤ��g�ǠP�W>���R�p��٬i�5HE��P3�!���W7f��7+�=�S�i.~�=�h���Y�я�t������m��L��:[� ^���U��S���w��C��#� ���&d�7.����I���
]���n�U�;
�R)��X�z�Oh*�d�J�~g�� c�FM��x�|/l�R���PK���I�H��=����I��8<� ��}*�Z�I�wI0�-۸�8l�兀ůͤ5�e+���I���D�g,�0�G�iK֡%��MםCy����GˢD;=J��o�1HYQL�����.�vT��bZ�L��5��
Hg$�I�}*�,������d� 