XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0?/��V��/� �ː,k�+�Lot�
NA֓&3�s��x����D���E�U��Ğ=�/6I�EB�K�u
Hb�I3�z[���r��L5����tz�|Wh�m�O9�YbA�P~	gfg�p��i$A�X|���j�Àr�sށ�s��K��-0`~;�]��$l6תk�p�b����CSL�MR�̠���&�IT�fM����݇��?y��8�(�\��\��:d�]�#���0 do-��ڠb6oO�cY	�.����Va5��Xm]�Jg@�� <c�� Ս�y+�K���Ix�,����I��B��` �D���1b���f����\[���Y�tMD�y�MP������$��JZ���k���ln�Ø;�2[��*�5AC���&��F��Tu˱"���Yh��]�2�!���J�ed�b�p8i��C9�U�Vo��|!0D��WwsG�>�Wq(%�O%.�Mf�Ѵ���������xrf.�_i%�]�fg�*y��:a;lڱ5���Z��ݨt 5^B�	�M"���o��5�#t�0��z��/�-�q�l&���j��$�2�w�5����ly���7|>�+EF2u;2w�[�w����'�eCf������Q��X<�x� 3P��l6�	��R���Й�ɡ���Q��FɫOV�����LD���h�K�hké��9C��zj�|5�4�3H��:4� �Q�1p�`�+a��m�`YU�F�K�������f�~�%jH��PԁR�XlxVHYEB     634     250@��v�&��^�,������
� �.�_�/wT�h��b�8��MH�S�#H]%�Pu~Nr�T�b#�����~*��]�N�.�ŋ v}��>v���2�	-0����6�6X&����|s*�-=��A�̲�<��χ1@��3@u����ӬQ�r�� �X�Q��ў�	5\	�(�+��c��P�e�Zɭm�hB�v�$@|�O��aWL^G}�O�ɀ�f�W{��F`�;~7���Y���u�P�	Q�Pdμwn�f i�ew�
S����� )�4R�ҩʨ���|uv��75 |pJ;M%X�GD)�Z�M"d��>��1Q`�Э,?MHF	�-ۂ�t;rC��ֶ�q���6K��� �lk�j(�R�8�������w2���b�̱*<��������rn��άB|��U�k['�3K���3��Ez����Y�x�	�Y�&Ko�����
d�xp�l���+	��в�d{�Br��}Xnd+�#,F*:���~r8��J�R��p����Js�Gп�ފ�T|\�[��_i\iU�����'��?����`�
�iK���i��L�