XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�?Cܽ��+�J+m���d4��{J���u�D�A��`��\�^e�~���Y�M!O��U�+�>[�O��
O��OǨT	]��:%��CoRȴ@uA.����8X�X�Ϭ5��6'���*��xj\�e x�B���7���1��z��i��ĉ�&Y�&�ܖ|2ӥ�^�a�H~~��=HhB'�䱟{��X����'HjQ�	�gez�;���;:n�{B����I%��x�4PLE5�?/�=o�]O�H�[R�
uN�ɫ�c&�FF�h�R�'�6�����]҇�З�{���=s^�]��~�9P�j��io�'"���~���Z�{j��m��4��<� 1I1=5՗�e���l���p��+�R���a�#�z#�B��ހC-�#Xa�OY�E��zz����\��F���.��5�Zzf��E>Hb@OF��9,�1�-&�y\@ ��I�c(���������di#q�qƸ�&�#)Ȧ�񠏪��φ�O安�M0����9VD/vi�,5��f߽�_9σ<��:m<`@��*ۧ�i�.��?�pNA��Ů����*��C�S�u�����Bw��
u�_v(��S~�lO��Ae��nM	o$�D#N�O���h�K	���ί�~ �itw��Q�$޹]�dD�g4�Sb�p{G��tt6�5O�mA��6����U���1�H7����ɹӦ�K\*ZF|�C��i%��7�F������ߊ˟�����Z�qw%�.>���^���XlxVHYEB    3a1c     d40Yd%,ytj.R$��c �t��-'ۗ6�Uy�Q4���ǕRoY�!�ĪU.ː�ͤi���퓮ֳ\��h�i�搻F�]�[+�Ui�J�_!�t�pn�М�Q�*:��^����e��!ǦUz������;�ux�|N�3�#��r�T)��"��2T��74�c�����r�w�M��
�1�ע����Z�=@�^��w]������,|Q����G����&t���,�H]�e���.PH��B�A��ǰ������JX� ͞`\|bU��,'w4Fͱ@Y�\��ٵT�m��ʡ
��b�uj���2n�V�Z&U �+���)IՇձ���0���	}K�������o�}N)�i&�R���`�ex�R80E�=ܣ{$��!�ێu�t�}��~��${�b��@`�>�K�#�� �Ƶs��,:��v����Ϟ�����X�s�C[n���3b�W�����RMbu� �9�	Q$��j�_�W��`o�
=}���H�z=�_�%��*(��k�5����</�u��@J�M����x�gA�26=�LeM��y��y#F}�� �'��������7Gl�"�q�a;K�,I�ˬ
�gv�� ��g�"�h���"]W�%;l�Ui�n%vD�y�Ѩ��-SՉ�� �ׄ�Q�T��U>H��j4d�ź4�30�<ܤ����4j��&3�[���Q��K"t�|#\, ��d�!&������y�`��q~�N���h)�I.l�<A�Yf�44���>[����A.)|Q-&S�R��86bSc+�b����2+:�m݅���*'9��٬�f)�.��s�{�P��|����r�`�3����k�.����ч��GԄ���j�KEF�ؽh/��V��;WdL�y),B��L��ش,r�-���O�(z�b��.С߀tjeD<��25�X���(桒���C��_���s�������!=@�l1����;��DD���om��P����U�Rz7/��`�ܩ������D���+��l8G�4'{�>���l!��m�j������8'(�D�7-Ů3�E���Ē�Y��K��b��pWM�!u��ț�K03��e�_za�y+��U&����=&���|Z�Hf��򦌲?,�NtW*-G�)����D!1�%���{D� ~+ؼ8u�#e� �?�^/��ЊN�>	*�V����x���z,��H�p��:����f�C�#dh�|j�נ7�{��r�I��3<$�H�ܶg�C}����:�%nj�冢Wg���.�=�4��x�\@��Q�T���*��xM�ĳ�ԯ���D��_@��D���I	F��T���A�h8�m�dId�H<md���.)����a�r*M�Lm���'�NbdhPg��ځv'���Nѹ~I~8'�Z,��-a��0 B�eh_����UUzcr0���ϘBK�%U�0s�>��Ei�o�s_j3�SĻ��ٱSj��E� �a1�Ko��^r��O���nS?� �]�-ybH�+I�	|���I����_jϵ�x���ζ�qe����o;�wI�n��8�v>�pǿu�O{+���D/�(M����O柤��+�^��| lE	U�Wl6?��I`e�@���@�u)��D�����-��Eg��ߜ�u� �q\k�&�P���,�ڲcK��#履��@���F,�.�k[���O>�08�c9�7C��N�vK��,
6����<����dZ�e�_e�^��I<�;���{���n�{���R���a��R�Ҩ�m�9.l4�~\�` �O�	u�z3>���?��k���+��^�tN�(!������d�!��l�Fg��b5�
�S����N%:�(4�!/j��d�I���l�.�$��"5�{�;@ς�C+}t��<�03)5�f���~�p�N���܉��`�[���J75�0��7���Wg���Ӫ�q����������\���)`n{�k-�æEIL/6�$�u5w���2�f�����h�/c���:�H���֑k��_���y�c��9��_�\��sԕ^a5�]Y��X�!���nhQEG[r�i*v�˼�z�r��׉�K�8��7��5���������y]�>�-��&Ӂ���P�4>R�0+�Ҥ��f�Ԅ����MO̘VTh���{1t�)Y�*w��U'(�3�?� M湲��1�B.d��)L��o���NI_����߉�0��bO3 ��*0��m�,��.j�5��m�@�Ghj�ޜ�5�YnC�8��HP{w�c����Gq�70���+"��jl��Ed��W�+=��X�L�N������,͂�-Z#�UF$����ez�ტ� �N ��5pQ@�Z��f�����T�b���H��87����@��ǚL���jv�-�3��r!N�£9�/�v�e�db��,��X�D~ߠ����&�aW�C���	a*W܆�!��8"�E�wn��~Ӿa��(�u��A[�¾MI��X��?�_;Pf;��U#i���YV.?�M]�q��o"_����jr�S�vD�R�o��s�N���Co�(<�#J�J���l]!Z�޹m��߱	-�dL����l��xq�r{dэ�UO����fJ�ξO��h��WϨ/���K�)wo4����n:z���,Q��V�冇0� @�����3����i�0� ����V�uG�P���&��޴|\龑@5-�UW�ɨ�m��\�9?]d��G�͵oP���ֹ���
�oT	|e�`���he)C䱱��C���gB��"�ng6��\���'Ps���[p�V٥�@�5H�YJ�_4AJ��5@��%�����ǯ\]Ξ�$�M�LJ���I^�l'"�J�s�Ps��=�&紸�U.C����<��k5~r���*Ι5#�[�\��� i|����M�(-��f<Q�`|�83���HI�i^�sƺ|bI�?zjv���~�5��n�:'�h��(+n��E �R�K�:Z}��>�k���^hC+6�CV����M4Y��|�k��f���_Oą�N�!�N^�~絡�w�%fH���\?ȗq��HY-I��Y��Gx���ă���:rӵ�����w��4��Y����ݼH�L����GW�5���̉r��������`/��q�7�����t�ܦ?�P�k�M�[���%C��c6�~%Q���Ů� 
���>�-\�ԃ��+���q0���	��hǫ%�L��ͰK�v��J����?�èj�U_1C�!�0��x�m:�l��M�A4k��,m4�o�����b�XO=��=O�?��?�H��s��"-�˘/