XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����k|��Q��Tb�y�_[Qy3`?�z�IK̺�l+N��m.y'q��n���C���]ڎ�
���C�np���#�?]�Q��'_0��By�5h�J�X�ǔ�R�GD@�6��{��:�7T�&+-��B���7d*D����k���L�v��̹�ܚy�s�� ���j�}�h�Xt�u��\���Ȓ��fE��<.�&�=�}� k�Lx�=�äj�B����D�6��]�ΑvN"��ia�`9Yn���I]�	�dO� �.�Q7�Pb"U��y���%Z�/�3�(�3���]ʙ̴lG=8�E`�i�Sd����0�&�.*�D "���� �vC�߈���������~����MR�[uP�5+<,(W�&N��2�!M����4kN8Q��s��瓄��:�귺���� �pM*�����o��5*���U�²���~)���e���6��R����E'�a��2����P��R�C-�-*�O���7���;�����t���..]�:Rg&/N�7@��w�>R�Y1EG[����Hi����a8R���/5$Rԟ>B�9�,�~hsN�o��v�|w�R�(ȘALxMշ�^�p��/)9h�&%ͧg99,k`��c�a壨`d�m$;���buSF^qd��9��y�Y����=�j��m��Q]��h�9�R��)���闳A�*�-	��I�=6�g>�Cy�����v�9t�㋷L��GO���YR+���Н�.X�ڂ�k����px�XlxVHYEB     a56     380�S��z�.Ax��[U���0�e�-�[q��#��o�V�E�r��y�9K0�Qb��|Π�V,$���U�A���4kt�gJq�}O#�N�(=�/ښcy�G���A��Kك���8"�%�qZ<a�����`]��_iL^����oq�����'zd�ǝ�CWN�0�d g�6�-�P��t�ʤm��	����t������%��jh�S4�+�@�oU>���{F�A0,��-ڬ7�"���ID�pK+�Nmz�v�ܮ����Qa����a5H�1�v,^�������`\�t�PFr�X�9p��������\�^E���m�D)�cׯ�.j���O4~�8��1ӠVl_ɀz#�I��ї�&"�{W�ْ��+� A����,>]��x	�S2/^�nE.Й��ͬ
�6�W_ό���4���l�#���p��B��\����vo��yZ][c��}GaL����=�|�Ze\50�THda@=�T{+�J �HH�>q���U�Sq�*�u�Q,�(Yy�,��x���A��\�B�9�Rݖp߼;��	W_>�b�%u,��� �pK�r�0�Ӟd ��vu�+'�H�.xݎ��ɹ��1"��Y{&����m�E���)H���%-���Kl�F�����嬵���k)�Wx)U���@ڪQ�F����S���5F:�bP�� ����ec��Խ]�p$�<��]7+�n)��o�x��BG@�&60��F.�$��5�L,��f��5$.���
�ф��������H3��ô-o�[nUm��$(~��>	 =G?rXY=�����B��M��^�4ޖ�h����@r�*�d���4��>+�]8Rn����f�����8k�>H�{�������^��ُ�֧H��y�X�Kq