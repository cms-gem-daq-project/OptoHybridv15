XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���aXݰ_��6�V{�uVO���Q�����7!h�G���<��U�V&¹��Q�3;U�^p}�4,��&F��U؆��6�H����\V��J����C&ֶ7��Q7�@8|
�PC��9+h�\�^d)'��E4K2sw�tw�r2�H��0
���T����$V��..��D.l����k3:Ѕ6F�I�ƴ8��YM��@*���q�.��j��^@�T;sU�G����B<��� �P�l��몌���;�F�<܇VO��w�c�ծ0�8fl�b�	R3���8v�����9P[����E���Ą��L'�Y��:G9~T� �y8�.H\�����i�L��xl�`BD,#xrj�fD����\;���J�
��o����jrvZn�+W�n�A&١6� ����D?��%7b�m���>k�z�f�՗��\	k����8b�q��?��Pv���K&wf�)1$�r��γ���t���}�=���+)���93��������� 6����%,B�q����U�A�u� �o�P�W�З:���-+��(-��Ԕ;-���d[�����ˉ˂8��}�2w%B5x�9���¸�=�kZ-L�P�'�=3m�v�*�E�,i��"�Ϛ��ǧP������2wg�JzA[u���-�A*�Xf��А%���3����|�
oNҝl�i�{M1��n&����$ټ�9��e8�ŷ����6�Oy>��ȥ��~
�
�!
+��e�V�����0XlxVHYEB    7e17     de0d�z]�߶ɩ��%��N�����g��o��%��
XҨj〈J��~UY�^�VFr�ilЪ���O�G/0X���8`ךmmw׈V�Cu*+���!e�ͱ��%1�S���v��T������^�#o�A%���&�qa� �����,K�7�Za`��\N�p�VqU���P��[D�����㜒0i�Q�@[�[䲮������/�
� e����G��݌XN'+
�"�u�7Fk�h�58;�BR���XŮ��~�[CS�t�]�¼��Md���wo��g sQ��>�@���}�1Pwr�����mz�f��2�'�
K�����������U�+^ !��=GtX�"����)�VJK�K�os�mI�d��]�&����Mx4����q��gʦW�e��H���r��Z!�����]|]��P�P�-��E'@���Zm�3ֽݴ����Jȕ���-B��&��[P��v��6O��l>Ƌ���7�J�zeGE搏�=�~�m���8o]s!*�r��d�ZG>�F�8�Rˀ��1�+ �|/ܽ`mܹ`%�v�K%t��ŀ�fӿ�
Fed[=[f��Knj<�6��ը�;6�>���ث���n��\{5!�"^��g�Lr�c�5�d�@DL4�(�\�w�?�7������Ť�IpH��0�����k�V�Z��TS�\@���2&��]3���۴�����*����yZ��!kkaǭ�Zrj��V1p�=N:��
�G�ݺ1/.����;[���e�����w�O��,J�%M5E��Q�m�Hĺ�0}��<=b��\���{v+�m�ِ��)ӳe�MYɼi=+ҟm�>SA��R���"��"Z�N��w�G+[�ˠ�ĳf�R�B�ҩ�EB=�GFY��! �4�o�r��j�-����w�å��-���+ �N[D{wgk1�p��$Al�!v~��ش���e�_�ttGI �3c[#q��Sle�6a����x6�a+��.E����w:�m"�r���i�Oi|L�=pH�]:���T#�b�� .b�2p�H�2f�Y�0�¿>�ѽ�c����_��L���t�9��b�2��E�4n��Z��T��l�2�u�P�C#h0V�5 ����*�}��"!GngRr�q@W(��i�rq�����H�8���hb-�?�^:��
�)k�&LqJs���#�� ո��� �'��O�S�'�$*�h����{��o`�36���+ڮ{�E\�$d����v�9_m��dK_� .wX���)��$|E���:�e��%e��D@��_�O��ܡH׷��}�ۘ���9�4Cq�5
��g-O�x1ٛ	0]~t�b/Ip�1~�Y�$x^#B)����Vͳ�}u}�5�2��y��Ŭb����,@E�)9 o���c3��l��5}^c���iS����/ӝ�[�fNݻm�d?"K��1�ƅٳ�G���i��2�N��w��ܢ�U�y1���)L��e�n���'B�mn��f��*�[����|�~4��L���A��/�0[?���~��2i���b�?�, eT���]�	��\��S�e�,p��=bBs�����uo`�dkq�,���~H�k�?R�	����_��)�z8��Bukh��Y?��L{ʵ�5���Z���'w�\$�'&q��WK�Y��&�2Z>��+⼝��E����2G�#rl�D۱p�r�%�/��<|F�;����w������F�y�^�e
���!�?�	�jY�6l�^VS���=���,����CG��Y�D��=&�V��ś�{��8d���3H>�1mI #�=�,1r�UV�\�3=���\��u�-4k�gT�č>A��hUܴ�� ��M��Dl9Ԭ3Y�����d���y��G�w���@zZ�<�p׾�x�|�,�x?,�[1��u(�9�,�����\5a>S��!��u�����|}7���e�*�t������� C��dT�:єA������/	 �D�+��`�M�<�1U!�"����������pG�/���,q�D��0XvQ�>EHL�L ั(��.��	��"�P�����T3K�\)�4���]0T��Ancx2�2� 41"C���1i�v�*��4�P�*/���*�YE�M�7\$|�J5�=���{ģ^Zd�11,�Q;��Mp1N�\$��d>0h0�f{���1Z��[q�g
Ъp�ԯ�����AU;w�/��:��
*M���>��*4�F ,l2>߯�"-�[�D��#��*�9�)���҈00��fL	��{e}�J�8���"
W9,� j��X%��qO�ڈ3�=�
��u(���5���Z�PI�m���\K���W��g��ѕ������.��(�>��[�\��7a�t���{�+���
��!;�iy�v�����.����jA���V���*Dq��2UWRn�sۥ�;���R#�L�V�g*/<���=�A��NM�#��+�P�f8��U��N�0
�C6Ks�p�ְ�w�Š��9�+(x�(���Ί�#G��@Iv��y�&'-	��`�7�TBz1�������z&���r�qδu��S3��=�FXX�L|uf�8��?6PCXy��븈R��nG~��B�j��4(8Z���xݵ	��a��y�$�[���@��!4$-�V�����c�<�����$��N��\Г����X*Q)�O[�ʞ�Nd�� R��z_��&�9hE\]=�P�Vp85�gK%�!맡����0��V�3��L��oM߫�����X���6�����j��&#�?h�9�f1��phT��_�N�z�9˦ky��ї���	��b�Ey%E�:��z�`d�-�2��}r&���
�X,�� �)��
!);�.oI~�9׋% w퉘�����
���G,�矙���G��sr�#:�Y�H�����Y�F��C�������Vm�`����֫�n>��`��Ab9�}�<�^K���P����x���YӖk�]���8%"���Y�t��+�b5҈�� }1�}^|���.�:ְ�s��-_[�}�6�#�,&b#�O8��KTi%q�3�� ,�J!r�
ĞC�-=�|w�+�����bM�׆�����P���n�I�����V��S�6�F|$�Q[g�K�h��s��#��)�����p  Y��oDPb���$��x�j�@�p�Uq#"yZ���\ϐ��qB���@3W�*d	��P2~
��E�?��w�ͽ��
	�5C��W5����G���$�3.:G�C�f�i4#h^.Jd��3-�[�	^�i5�Y���ӳRM���tc�Ux��1�H�D����W)���#��� �l��o�E@�Viݿ����~Q?��2����T'�7�dթ��!iŽ	�fY���Z6G�rkAv�2}@F�iQ$�)���i�����mw�a1�'Hw啥�J-W���