XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s���*�����}`�A�w�[�SNR��U���!=�I�l���J��̎���d�qꈂ��ƛ���T�3=/)K֢�&g9˽>��R�!�w9�# �I�Bs3��Nb��x�24�P�!��	U�>�4S�p�Θ� Q���q@�r|�ane/�r�X���Z�*�gv�e\���}G>���ٽ��P��/Ũ�{Ĳ��(�D��Z*�̽B)-%�Ȼ���'�?�ț;}��T���_DH��/�p����E� ��Wh�f�yS�A�&��.����XԆt�$��	w�X�ˆI��������#��W6��n�R�J�ظneK-�o�E�EHi;�OPٻF�� ���-tcN��5;u��kj��3�8F�.�Fp!��kPs)��ʃ��U4�\����ǥD�kez��Ib�F�-��ʌ���R'A4t�;+gFN[!I����2�%�oݖﺯ�}P�E0B�2<�d��� �P�G��n�ͱǲ���t�Zݰe=��傉t�(��g"L�GPߐ2�˶MỦ���[\����o��J�H),r@�#~�M�����SY��Ep��(�1������������c<'&�rb4�}Ԫ�vִ�N�M�{4p��e��-�N��UF��f���z����h��H�I+]38�[6Xi�����; �Ƽ�״˶��a�LC=Z���L�#?s��Y۾��U�x=����%{|;'���%�7f� Q���ő���)��yQXlxVHYEB    b892    1b20�	��3��'�f��f��p�8j��H�~��p�߇��ܬ��H�b����j���	'�e�~���XP�d� ���N��4����ˀ�0A�q��.�S|��.z1�$�'��x'L�����N��]T����[��d�84�~D��:���Y��wx+Ǒ{N{%i��A�w�մ=Ά��t��Z�����l�Q ��)������������S�;�1ZG��;aD��e$ �>#�K ^��Vt9�,?#����;x���4�UA�����#M7-�Z�Q�E����
'�E�X�3!�|[��q��菩�Id�2i��F@���{+6�P>}R[���.��Tツv8��ɡ�v���N�W�9b�F0Ɉ%d| �����7�hg��{�yol�?�*��6���C��/��i�]�ʅO��Q�vX
��?Wg^;�q44Q�F���_�eh=H��QR���"�D(�k�h~AL:��ʜ�bPN�",�������(@��FOq��I2ٽ?�ix��#O3�c�T�^V�o�k�OD|�X�Z�w��'5�'����˥�b����y�j�OOiSx�.-7�,��@-cpip��N"�Ms;��@���@|"j٧� C����t��Esb�(�M�Yt���Ar�f�ԃ��2=K���^,���&,� p��'��c�$δ��a~/�"a���2�#�����! F h��V��B%x�
?|k��U�~�����2E`uP\�t�H����]�;9$rn��ؔ�h����̱�a^��G/n!"/��op�b}�U����������Vfzq>�����3F.��e�̈��A=PkV?�@9�J,4X�}�q�4�.cZ�|��`�f���4!?ܯ�y�} %�;~9� ~c��m���O�%�����!E�,�d�?T�C")��-�, ��]h�dN�~�(�09� o�FH�+�EV���D��V����pS�`k���������#�MW��sFn����=����4�"�c`�E�����Ca��yo��A5=2�B~�$m���i�R�U8C�$^��T�V���<W��gc0�wܶs���n�jr.QyGt+�u �Ӵ�Ć:/�BN	��=�S�Rs~��V��N)è?U腰���@FQX���v��\�������l�J���¶(����@WX�G���t#x�]V��-!��T���H��N�3�ݸ�h��ػ��l��je@�w��t��(jO<�of�ƶ'��o�V���Y�`�YtY8bh�&��rC����|4r���F3>c���ZV�??H�(&7e��G���;���~��~L����\��ƭm]�쪾�C+U������ ?�9��Е�G�%ui��S�qo|��	KΒ3M��n�ϒ��M�(>	b�2D�$E#NFiP�p����2U;k�W 2~(���z�:%���U��"�,���9�J:�����T�P :��r�	���ݐ��	�}1�hߑ��4 �U��<D�?|��
��
�yҌU��'����k�x���)�"�	e���z^yv�-=�>���g<E�>fo�Gfx�Mr�FY��G���UӜ���`���v�$.h=�?M�ܢ,�"q��]^��V�&Q��O<ĝ����X}���Əs�%��3dN�i��{��"�Q�NP�a�o�B�R�GT�)R�[
�?��unf2T�>H���x�]�U��BUo�!C�ƶ��]���గ���#� �{/�&�/�L�M���Ű�wg{�����v�#���?�'���M%�w@d��A��i��o����YD3iZ��$�UC���m�$n �X.y��k;�Q+Zi澋�<��gu��4�j6mOS��@��%u��3�MM�g��U���+Ɨ�|�rV2b�����hG��T�Ơ���F����wm�mpC7�a��Ɖ�y��q��m9kU;9�xX4Hi)��qG��?��hs�]�#������$S�(}�����]�m�Zh���R(�a���/;�혘�6�p?0`=P1��y}�mC�"�B��u�h�,�v ��Y��^eK�m����j���z��]�L��z@R�-����2za�8�B�^�屫�(�{X�5�	[�-���^R$~aj�U`x��_�*��]���Ej�'�3�'�V�+��(�Ce��\����a�y���n�K��מ�q&�-��Yw����:>����*��ܲ�����e�-ʕ�������j�����ݩ���|���(g���B�%�Ȩ�I_���Fd���v��~�WL��V�I���C)鶾��:Vk���%lhBL/���>�̈�Q	lF~��Ґ������ǽaf.(*���X�_C#���i�i����f�JW�ճ�&�"KJo�s۟�č��#��ڱTe����ϋظG!��"o���詫�De���fh�<C�MM_ڸ����j�e�һkk��<L�D�))��NCڌ"lzS�8��ښY�p�P�X�ޞ�o5��V�
���c.A2��/���݆m)تMP�����|{~��"����j8�����m��5���x>��3��0G�<��ǝ�*v��s��sq#ݥ�)�I�I��֬����l�!�6})��m��Ao�J�N��J���S�Ꞧ�f(���R\d���b�o�TcnY�'����s`.3BǾ��^�/�L,ϖ�.Y�i9&͛}�vK��4�Q}�����\g�0��&n�*�<�elr�-�lc��9
�e�2i�8�U
���׆�ܪ�eS$�~�*L�D�A��l����t��&��vD��JPE����M���RױA������0N+��~BǌI ��̌���\\�����p��&�ly<u���i�i�{dy]� ċ���ݴRG\�IQ�?�>2��|�:ڍs��4\ZҮ�@_��������L���Z�)���$^9�wn�DAW��:�"sR>%h���x����JEJ��Ҝ�U��ߩ�6FvG�� Pe�_$��ֿ�3���b%Z�ޔ��yW��l��z�%��=G5�X	�"m�K�w i;y)9n��Yp�)A/�6������}p%E�:7����aݢp��%�]=�VWr���1�`~��/��{��	C�Ž�Oc�W>u��g
��d�3���Ӱ�umRh#�<ɺ�؈��BE��,NT]��xbS1G�"%ɈU���T#�`�k)�4dתj���@�7C�O�OñR>G]Ꜽ�G��N�<S
���$���/�2#A�{|��+\+������I����>k%
6�Քc�x|�'"y������i�CWs�г�]� o��+�����[SR�Ǝ�N�%��b�������ѡ6/簦��4ϥrTF�հ��Xг�D�����BE�<</��H�P���T�$�F�\gR�TsE�W��GM�X"l(޿x*��2�ק�~�.	�ڌ0w��ێҟ��5?��)U�(X�W���jPӤ�^��9�kl�L�|��4�ʼ*���o@��~UJ&�\v�mF�-p�9)f~A��QE��P
 0n��ܒ/�	ֻ���%ʃ,o����~_v˲q<��ҸC�z탢i�q�8{�o����|2�l#wp&OS��Q��o����/4�M�ԧ�ŀ�!��ni,e�K{~T!�߷�Y����/��od6	Ao>�`��5���͞�9�):�:�e��	�����s�u 'עB�l�SL��ˍ�}���vI��Ȼ��Z���6�#����U���?�,����nc��ՇX�H9�Â����k^���[�T����Z����Px�^�O���ӎ�+Ļ���i���E�:�X?�2��?h۔��WN�390���v����U�o�xK�Qjb�ڡ�^5Ll���󁽠d��r#�k��5��bJG���Xe�XEB���0R�h?�Zbi�Ru껅˅L���Jf~Af����h���-R@���/��S���2<g~Bo�.��V@����.�xuuΥu
���Ѯڦ��"@u� {�dF�Fp�^�ȑ�����1���SJ�o�fS�JE`~:���$�O�U�\��}���mLJ��t�/�i��6t�� �^���f;�a�)ŀ+��%r����������*���e���;v���'cq
-���� L�ۢ��p%5G�S�	v¿'jB��Y�R��#��a�.��o�g�F�������ldX=���r,�t��|)U�(��JA�S�6����qg����û�� ҵW�>C�> 6�_�*>%Z�U�yO�9��f�����S0���*�������0���~�4
aj<Y�.c�3)�����'�$����� ��֋��f�F���V�s��Oү�v���0J���]�"�B�Yp��QkO���=
�%�g�c6�>�h��?���8�R��������M��{�Ó�O�$��RKD0L��zf��3S�Q*Տ���"הϰ�e��O�/"t�ӱ�D�$äf׽�`e��$���P)y�/�f����<7T¾�e��S.�9��}���}��/%���Z^����_���@y����K<ŗZ)�T#�{EN��)J�jYZ����
�~X�"���m��]X~��w+)0�}�W /�	ߒ�����G��k��s�k�Z9��4BkҞۗ�M�_��	�Ԅ d�?,}<��F��jf�?���H\>�0P���<��u2�7����[O�M�X������� ��Ss��z�-�SOw0g� �Q�S�A���i�$k����DbhlRh�̗#���XGә��d�hɸj�M��'�[�K��l=<A���ڬ�����}�t<�{�E=��e�Z03�iٵpK�	7n�3�"q�����l�N���E,f%��Ɗ��p6�h�:�P"0�f�#����7�zG16�NH��TAfi�A�8�˘��i^U��F.������@��E!�Q���S��1���A6J�ܓC_׺�H���=�U}[`&l�I&C��2�v�a�>�����8o-<��Le���#THߜ�+��Iν��!��{��w=�;o�^'�0j�MV9�M"�p��`���\1�g5��Xj����썥]�H�qf@��&��M�����	�6,r\,�^��mA��Y#�:F�B����Z����x- ��ܙF3}��	���C�n�$�K;�j�W�L������	S�C(�6���i������JS����fuQ�S�*�����Z0L��eʾ�ȝQ�@��D�-]Q�%���M��v��S�������+M���U�v�	(���������!ԨJ�� Aۮ<�Mrm2�̕�@Òـ�OT������K
G61�ox A�A[�.N r��ĝ�>#D�jsR����p^ώ�����ѱ��_;��+���j��4)g4Oϖ�)U`9�|�?�v���\�4~*UL/h�B*��4�m��M�r9�Qf�tG��E'ﴮ�eG����#t�� .� �t
!W!\���NQ�Ψ�c2gJ��d�zͽ�2}¶�f-�?�`$'��.ʌ�2^�{\K��^1�����є+�uf��J�m@)�����������>h��E-F��s��鈃����!�f�bƳa��s 4���6/��+�?)�DFZ���@�l{��h�%��a�J7(˵Ym��"��ʁʣ;���4̹j�Z�ljS<\�J*,���6���>��uDP�����@�)�����i�������H �08�Y$�-ף�[x��ɐ��>������6�$%���ayy�`��r��cc�j6�DE��p�_�w5Zs������N���a8I��9F�ZU���O�05��Q~�<]��h}٢P��Y}��P[���s��cPR��N����5�b�줐�Ř���3����C�-���[5A>�S��.��(4G�n���R4�4Q����0̒�5����R$����@�yu�7q���,e|M|�i�yi}�B��q��������(���7�UN� Pԙ�3���/tM))�Z��W@�C���S�N<I�Zq;�m��^Os
����b˰ǳy�Ð���&#�/�#�נF������x��{ۢ3�T?�_��M���aLQ�_y���fy���d֋��G�V�H�W�M�Gw9�s����`�I8�T�2���vkN'�����8� io�wҟ�m��G���z����P�B�zP4���j��C�ݜ�OkЀxU�j�.A�_U�{f� �9F�߇g�e��Ȫ��R�i��P�$`�!�E���-��mr��w]��f�[�HF���d��,ʪ�#OTĲ�\J)�WR�|x`hA���,J0�	@��DY^.62묀�>6y�����l�ޡtV���S���b�q,�}:G
t��5�IQϯuQ5��J����m~��͡(k>�B҉��y�5w1j���fu�ԟ�*�������3+��=�P�@6����H�V'e�>o���+�M�d!��A��^�I��gs|W-��E�|���KoH�:�wZM��äp�%�$��R\�&��a+��c*w;G^C���tp*}����F�Q���Qڙ2B|2�6�L)���g�x=�������<=�Q{�Q����%��;���wɺt��0N�]��6^�[>=5�+���I���rt蝙����<�<�M�����[t5�j�N��z�j���I��Χ��j�v�r�Ƿ���d�#2��Xsr���78�A�M~oT��zT���
�*^?y�V�T����%o�ɍm.Pq_��1�;���WgOf�=�TM
��M�֭TX����Q��VK��X3fn��Oh�h�2��^��k�?�KR�A;ʗ�p�