XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3��������V"?�FLqe�N�Ý��H���;HY�}��g�V���v>�6�-'�_��P�5J�"��k�Z�����+ho Ma��$םf�'�T ��E���-���������Enk=���jc<����Cf��N���麈�v[Nvy,�@��{0|S��n�NA�e�o�e��q�x1r�B\tC��cyjG�<�n��|?C�m�Z��]U�G�t�lc�>S�rr�0�YČcH��Y^cJ��������k�-^Mʂ2��M���׃q�9�Vv��k��K;�_ೄA�Q�i�����dhuϻ�f�^��	YBٺ'Y�A �����ۧyy��`S�(���k���f}�X�#�}�|�v~���v���m�S���ѡƑ8����
�s��"L�j��$F�J���\�u6=�i�-�������W�\_�*�����#���/��K�_$�Ŀ�Ę!���
����Cri%X$+f�:�U�Z�h������]=m8-9+B	O��l�UrwP���'8Y�^�){��>F	�9����)�D���h�(`��7���?�f�ɵ#4��	z���v~��B޹mX�'Qow��Y��ZO�t1�Tt6�ĸ�Cq�1,j��[RK�[v(�aϽ�ՠ
2_D'�8��|=0�g/��ix��GhAP�x�'��iFj|��x�LM���k��5냱<M���+���g~;�+�0ĶE�16G�$h�Z!�6\Z�ʲu�pJW������$�b��V��?��߾y%���(:�+L+��MXlxVHYEB    5ff3    1040��3���KRd�ȗO+te�
ӾH3_쵗A)��K���*G/�ue�/�-ޝ�T��.9����יOe��G�jjYQA;[�dTm6ڊ�ie13��U���e:0ή�}z6J���#(&������gM�{���¼�B���q����<�]�[����F!v�ߐ��������\_� A�(�p	���fד|!5)��C�h���,�TO����Bnف|B�v�M�=���3ݏC|.=�E� �[Ҋ>5~����K�~m#!-.��_*)�����sǏEx��;�I�E�Q[���ѯ�82�ǳ�5�Q�:/��j��ω	Յ���_������6��y<�Ǎ|E�i��m�����V�Z`��� p/SY;������|�J����url�77[���2^��ۚ2"��T��|�%�=�����q�m�rX��P��a�k�2�����,0j�p�;>��7�ӑ�!�--�$�R>�܂���S�Z�σ?�������f�aJ	���[Gr_8��=.1��iL�ɽx\�ڑ<0g�S�G	��I�h�:|+�b�Mo�N/?i�+�8c��M��Q�~xǬW�4Ia|�V�Z\������v:oZ��^B@3���WyA�u?�*�q� ���-�����ݨ��':��^%�P�Whg/��vixŵ}���"�w�S&7�[�j�OX�P^��L�bk_�GDR��:<�i�R9��b�W�����vv��J�]�f/��kcր��*���Q����V��_��L�M&��
fǘ�fɮE�jL�ӥ۬c�3N�(|Q.G�!�fY��;أ��nѦ��P�K5��CS�=n�m`ʠ�������Ȓ���y���I�khU@��4/��u�.1�����zއ.��Iۂ񣂴$ץ����4Cgpʃ������3bK�Pȋy����~�"&CK�[� �T�pE� A}m��!������H�{�0lͣ��!���Q�1�jUQ�A���A�ML�����g3���\�'ƻ#Au��//��udm���!��jx-�I�t_��.��X�t��$����g,���p�W�H�>AAV	k�ȼ�	�Cwm�"\��c�Y|ߩ�(��W�oT�بe�8N+�`���p�`!��Y���� !3+)H�i`��h�)%B����su�ə�χ�(�w�39�u���3Q8�%���������ǟj���:����\�{�ٸ�г\3'�C��nf�J�iͶ{Ў�q��qdI�z�<5nslծJ�M�N����wz{�}��MC4��=`�"��V'�|�	<�R.�cwo] ����"��f�$���!=hMϴ���X��#��'-�%�����o�7Mn�V�1��Ku;�E����
�Y�jIl�Q�q����Z(�NtG�('�7h���~���A��ɣ`�t"p�(WA�fm\��hx4
x�H=�m�,**/�;����#Tp��M�I�koD�.b����m�B�;O�<�
��{|���9.�]`��*��� ��y����*������Sd��<ʿ��j�VT�(#?�~�D'��w����oDv,�L�w��Q�� �^���������Q��������3��Jxjʹi��Tl���UM���]�޲7�L��}N�P||�ʣ��!�*I�S�t��Y�kYE��_��)I�6>/���Y���$�o�M�%��*���Շ���<p�׈�Ҍ��6�s��Єb��w�;���剌o�,�
4�������,����� �, 3�p�$B9�<�����Z��s
��g�\�|���k/��1�G�§J� 厩Q��
���1�8���x��Q�5nr�uPa��T�nM�0%kS6���lٷ�K\A�H�g�|ؑ��m�뤶+7�J�J)5'ۆXS�&�Z
�$b �f���q�.>��p�9_dӂW�6;���Ph�����yo���X����Ի�G�����n1��(�39��˗TQX��*ً��md�(�8��s�3�������g�PW� ֳ�%�6DC�_�
�ɒ	j� 1Qf��u�l�:I ��ݚ����FM����Z:
�q ����g��`��p�hgQ�ze���>[��
���Q�||�^�~4�[��jA�Q���w��9m�Y6����}��<�w��z�;��Ύ�C9���]�*�>�Hd�6to<�E�N��W�Ժ�Ο���4�\6���}У�ܩj4��wDpa
:�S��f�s!��A���FQ�� ��!�)�f�4��t���n�|!��<���XN�!S�������Z�rc�1��b��ߔ��$@_�K�ə�w�Mm�F���0��O�a��x��W��?�0���EQ��fL7PC�;<p � ���aUvK����WT��:��* ����70�"">��ȴ��m��`�r&�eX���K�(L�C[`���i{��XXUvJqv��`3�1���pm��mH:�>���nR���Yi�H��4u�m�Jo�#���{l\��yC-�N����٨�H�d�K�|s�ۅFM��g9K����?U�8�R�1�s�CܭF�9�S������	�l\_��뚫m2 -W�҅�Є{�J5��(����\�,���l\]��/���g���E.� ��m��p�!~O�.,�E,����-&�Z���ј4u��{�DM7�t$*H�n}������tR��Z�AՊ&�H<���!1/��Z��?�$x��u~=}��5��� �Ϣ9���:6�����Z#ӈ�<B�*�{���#]�pU�)� jg>��u��E�:j��VB�����x��pD����
�}a�������SB��NK`�!�MqPka�z��(��Du`�㜔�S�����vu3�4��s�%���|�`懬��,�A�.���bgv��0���Vy_��M���p�9���i���j~^�+#_3��қh����y��Z��
P6�fW�	���/�O�k�X4��<�����D�3ϲ�9�H�L�z�eV �rg��>w_�4~��� �Gi;�j���Ԑ��{<�Vh�zT���t��2��l�CP^�^��"N����
��e�6�a%�a���;�fu�S�����j�hH���P�Nڋ8qd��cHk�+l�S�.!Q
Z�m�g64}7efKg�|�:n<�������/6��N	�6N�$���x�����B�w���c�#�c��=iH��o���E�U_Y|$�5|{��r���d:��F�SfqJ��<"d�Fm��������Oy�T�&I�uy��M0��]���Y�P�!�]��& g�l6�[0�V�+*K�DH����w ���.����cM����	�?�χ&�㾿�����͉�m.*ʊ!�7]?���A��r鶢�E� uo|��z��Eʁ����L�Roe�3��P��V�n�R�8�C�!wv�_K!� ��G��;��&��tbn�V�`;TuŇ�9����hr��+��-t�|����CP���ɗ?Ѩ(��n�D��IN�y��h1' �m-������E�R��>��7�����d��Uy���M}�z�Di��ORl�,<L�wab��'�X�j
n���p�����/�/�������ֿ�	'��;���w�L�Ba9�I�צ�-ę�����֞|#������v�����XP�)�S
/�!�7���Wk�P90�i�����Ɇ�
g��p�~]L�&xL/U0FyT���Y�t� bΰ��v��G����X!/�m��6双-���&X��r6R��+���`�FJ��6��o���]`_6�K�NMJ�|����iw{��	��'���|�� :g��c�;�y'b�&��tu3��<;�>jP[� 	ʮ-�"��l���z��k�N�Ӣ��ҏ���4��ht�1����J���`xf��,w��EL����>	�Kl|
�4���]���g5")�Y��A?��5�&�IC����h>���N��L��'�F8d�ЊB�W�\4F���u��U3o���	nQG�=W�z8_�/�?�/s��^Y�jG��w�㳨M1Ō���2����