XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���l��@J��Q����Ff���A�ʛ�P�;1ܢi�=�JG��gh�j�n��:S��t,�����Pk=h�J�D��Z'e��{2QY�g[we�CR��� �Ģ\eŒ9	ș�&�7��� �ER�Ġ�E	��=#�̴V�`��^ϸ^���M�R�����ʰ��ą�*T� )"�����@��o ˀA��^�8�P6�ɰmMNm|R�|��Ѷ�[�5��<sm�Bۨ_侶���^cyb��il�+*�_4�gJ� 6�Ӆjk�W����Fu(נ*�XI/-���^�ȃcXd���J�b+��p}��Ll8h�Z��;R7nB������?o-���u�����؅��Է!C�����������>\��	M�K@��R0�3=e���H*)г����BQ�%ߋ���Ϡ`#�!��<y�:����`�-ġ]	=��X��e %��L��h3��OkH؜�����8�m��nH>�dJ�k��7_Ɂ���Y,���f��e�	v�3J2���a���4{�ik��w��O]5 *}J�Ƥ	4�����jB)[�z6�DT����S��IZ�@|�
�8�2��)�Y��{�s������tzS��.��U���o���%Ѣ�G�q��>���
�~򘬛� Q�騱��q�Z@��vnZfsd;��_4K�~���~��[f����#)��E⏖��~6�Fü�+٧�@�'n���@o�3���G��|�};_���XlxVHYEB    10ff     490!3L�=�E��K�۟Y��@��mw���s���l���(�uم�8�l�M�1��o�,۵`�����Bc#b͚p��x��>���yl�׌������4۟QH�DH�g[�n�{q���~�.7�9���W�񁙮8�Rqȋ����N뾒��U�V���V������p�w%˺z����m�8���M:�	$�۹�H��!�B��|��>�<��H�Ax�Ǝ'Js��b�}��~q'��I�t���d9<�;G6�}�˼=��_������e�����>w ���'G�# �3���j�(T0W�����x
��Oe�-6u�5⯷����.mu�Q��۴Cz����$�3yj�Ӈ+���Ј���P�B�-Jx�D��b�o�D��Q>@��z ҽA�1Q����3B�i��"i��i��Z�	��IC�p׾��q�hѯ�X8AW�;j��2�]�',x�nN�{D�x��`���[�"M��L����2�	�!��im������t�`)�����v�|��I,_�e�>����8�
5��TN5�'��9	aO��kD��֞�=��sq��r�Bf*B�m�NW�X����R8_4��U�ع�s-9��]L����>7��`Ï����
)�v>���&�b��e ���Y��3*�r��K_� ���w�X~��_�+����#S>hJ�����rKY&�ԸRY��9��U�g�t�7� 0�`��2���K[`*?9S>KH�`�E'���Q�Sz;��
"K+��gl�A�&��;�b8i>�0�^�s*(z⤸�P"h�*�.� �49�5��[��������xe~�*
�ާ��YTZ},��}k���?ЉK��^����"�A���B�����a���-e�A��wv��~���<2â�1�ܟ������Ne#-��3TF�[�_E��,��`��u�4���D	�;�A�V�n�B5�KA��
���^ion	T5��6���!�8K��?��B�(W]��CI5I28�H�1�	��BhPI�)�#E2R-51�c��3��8���VҌ�X�A /A�@�Y��d��iZ���N�S7��
Lt +|]����"�%x��ٔ�'��fzM���*��k������)jfm�-�����ְ.���'������;Ab
g�