XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ԯ�^�sq�昻��O:�����ȥhŕ�(c�b@�p�8�Lw����AWb?$74�9rTg����X��0�0-��ɏ 5���9X�D���KBvIK����=�u\�m9��ڼ�T*"M��3�8��� 8��>��;f.��L�!�/^��&����={|��8;P�yk>T��YD��x���eZ�TPp�M��~�	xso��X��,�U�&wh����c�����e����yl����K9 ��"$jF���@I�qb���#��}������Fjw�U���WP5q�f��N�o1X��E�t����
w,��ƴ))*Ѱ�Hx��d��7��I��� ���ꟺ�2΃q,�~k��q�y�;�k�L�{0xEw-�n��|�!e(�?��A�f�_~%ܲ��²��w6ޝY�$bJ�v?���e�/�H��;?�e����&Dsna�U�-��e�/�[�5�0lߦ����r��W��ga%c���{��r]���e�X�\ӑ�����H�"�2q���]p�@5ċ��D�s~;�E#b�B��I�%�o��`��A��"k���ӕ����-���t�RD�4yU6��΀�B�uhj����Ͱ��Ł#G�]�Y�e;�2����>��,t��to�����	������Y,
�5�������1C�g�h����;���!���&���H�Ќ�eC]"�S,�2�'b��LvO���N�B�@�?ј���J��ﷸ�"XlxVHYEB    1044     4a0���Plf���h�g����U�@�8P�����:#�ًk�;��_�Ȃ?�*<UŽܖRi�)�����o��5KȆ��M
fZX�^B�kH5
�n���s੝SC��	��a���XD�'�V�먜��SW��Y�����+\�ej<��羈���(�V!wΰ�yM�����(�!E|�PC��Pv~aؠ�	n�-��r6��P�忮{s�De{�ڝ�,���8i��5�̌3�0�O姀�gT�7�����2���b2� �u�P.����]]؆��S���e��W���f������@f���.�_��zK�sw#�]7P	�w�4x�v9���* ��o���n#���1��8N�-M �a#��aG)�v�.Py#r�2���z$]�_��B�`�	M�eX4����5��j{4ĵk���W�����#q7Or	< t	=��8����a�[��s�:�]H���������ߔ�v�1�,A��On��6T�,��S�bY\�3�w�b'B�x�~-+��x>�x�����@N墊�i�BݢV1D�ϭո��ݱ.�c��Tt=�,�zp~��J������o��D�Q�H�i���ʥn+*8X皲�3M��ž���M1>��H���Ԣ�����V(�</0���0�OI9{�c��r�^5��9���1��P��	
�I�(s9�؛�؅@&��ᄺ�V���4��	�ʯ�:���N�S�SvNE�	Pܖ;���+���ܷ�Qe�c��G���[q�<%��ϟgi��zs�<�<͹�ώ�'U�f�B1X����3&8)#������-h�l�x�Wn��i�*5�B��+4m9�A��#��7P�|��_*!��3xOE���A&�Z����e��@���z���X��;����Ę����$�,�����c����:m܁�i�s�\�L�x�޲!`��'�9&�m�<�Kт�W�(��j���5A^Ք�$.--b\�Ls	Ղ�j�}�`��)A�O#�E'����/�"�ه*<#~�X��^x�����G�M�`k�� ��V�w�.������A{��`Dײ�/H6�b������J�3x��<ͬ7�F"��kb�+,�a=g1*�� AjK�B���_�O�Գ���a�5;�)/� �