XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
5�,��Ӎɠ�CR�?	n�}>9 ��4Ӑ������A) eB��.9�m:*�,sw$�)ތ��\^�\��Y3�p'=1W�ys�Q�@7����A�.�k�9qp~�R�h�)��5#_Fv<J��i��)T�WfTf5����o7�u�9���f� ђX:��q�^[l�zH��I1�l`kA�e���)����](��P><�SZ����^U�W�-���#�Շ�cJ��_��Ek��d2Q��b����q;�T���.��_��o�P��7�Qj~N�:̹5��:=� �� 
��H���#kd�@�~��'>	D"�yK(f��7�mu��wX!<�O��+��Z�a�m�lz�ɽ�	65�KT�5!�+l68Lt\fb��t���O�͢*�e�{�\�wp�y^
�+k��SZM����M
.Pw�C�� ��s�:%����WE��|�p�A���?~t,����Vky{������|φ��?����&Nm�#`�.�����%��H�r����(�)y���aoA"�A6<�V�5���5���I�Q��U_��q�Sο�9��S��_�������d�g���1��8��TA3���$�,4�y����Yz�8��ị�>�R�-�ː���I54�51����H8bV^x��ϪGa=Q\-u_)`5�G�@�Q郧(��9iE5{Z�HB�/��	���	f�bĖ_�t4���}qR��t0����6L�RR麇�f��90!�'8�fK/\M_SGٴL�����ͮ�ؕXlxVHYEB    fa00    1a50l���d�s���T'�"�� �{�F�1c�����{��SI>|��j�:|}�~Ȭx�j5B���G�*`�T�V���F�joV6������El�9HGa���v?V��O�w�y�Ԫ�6HB.��B�������c�o����B�g&ԉ����"!"g3%�Ȕ�ܸ��9;g�{D��wM����.'D���w4������ ��}M6�<0��>�}Xև5�ֽf��V�"�*�d�ro��V�Ux����km��V�Gh�1j�=�E/��Y�p=��8+tbMC��E�*4�̪�vi5�g��0ǣ��J҉�K;��ZkFE�*|]��G�>vH����e��,O��]��D�u6-~R%���{�}b=�Q}�_�7�N�[�������1��C3_u�Z�8eJ���	��t��d��Q0'��ܝ*�l��2U�S�9�~"DhL�nϞ��Ѱy~�7%�c��q'�8DBl�.�8!.Q.��4"j�~b,��e��!��:�̹`���<f�9̿8����?F�!�HUub�>� ^z~�OQ�\�f�;���d�
���)h��~6�1�0 �H9�����L��p��uh�?���5
���X=h���E;��x������Q�]��g��!�[Y�ŕ�;%r��"�Э�I�{�FY4���9��2��ơ���sWnt�6�U���}��3#m�2�@�;VdR#�L��tL*JG4��\E�=L4@v��S��B<ʪ$��w�BN����q�F]n&-�`Ê��N퉧��F���!��ڥPC^[��ñA���%����_�b!x�x����2\��=�!��P����+3j!e��{��UU�VN,�&RN����A(�!k2'���j�X`�ÝJ�(uz^��ӊ-nW�.ۻ���><��쾬ך�|L��2g#�
0iC�K8��L#�)R�)<��򤢸ڲ@PzR}s��Ҫ~M�Ru5���x9mOgt�K�X��#�mb��<u��4��;�q�i)�f��ea�{��`!�����g��I�8�52�w��º�6�9��A%1;daL���0Q�)21�U�1�|$�U/N��yi��
]�p9.�
kNh.��C���$)]��O�l��&¾S��1�F�G��wM����H����P�9q6�~��������A=\5N�rb�a��4M�!u��� � ����'��F��3�
�@�,M��ꅡN��F�������"x��5G7�K�F/�����o����c�oó���+��G��,k?�nY��\�3	m6�!׆.P-���Kc�X2��q�q2	en��E��0�⁵��$��c�E��m�`m2�I���!%lH����dhj8)�_�{�|l�@=�����m+Nރ���ĝ�N3~'�2{,>�ץ��n���E�v�Dw	�T,��j�c�i~5�嗜�o�އ�	g�T��ۥ��v���#f�0cR �X��s�5���6�n^��g��_�0X~�>-��ߗ5�Ɛi��98�_t8���J/��@��Kڈ�P�
�#����r�Ւ
�c����ٗFM�jI�[yLk7
�R7cQLF�H�e��aG%m�X���	����F�-$�C>��@+׸�t"J���+KfS��#���� q��xoPM���V�<����
�H?v�S�8��/b"�[�x}ܢ㡐4�@� 准�<���znw���i}4H��V�b���{�m�����EI��[�Ϲ�˩Ľ�R�=�j
���\��B�:Z�$���x�Ir�P�v�3�L&��#{�����y�xGv#���:k"�2��N��}xSr�Y0�w(�K22��K+���Rƶ�:C+E?�>��7#"��ˏ�g�P����.9|,|!��V�^<��<��I��jV�*������94�>V)��}1��ITf�	���ͩ�����5�V��8�H[Ɨi �o���>����x.����b��Xh����RnRY����2v_t]�3a׍n+�'언���� 2~�(ϴ3�~y�t\ر���U��ݰ6>�Na�ª�R���	k�J�R1����:t���X��D4o~2��D�n4�ɿ�ꃪ��q�Zͷ%'���v���7�b=~z�� ��2��:2|D��V�Zh�4��^��W%�
��X����f�0��<R;���=�� oq�[4B=kp=�7a��1��|+��\��%� /P��2�j� d��I���7��Ac�2�+b��/�\�{�b}K���_HP�1_�a�N��J���An/=3��Y�oG�����jͯi��a����; �\a�?����A`[#���z1Zig	�<�����
���B!wVH_�<�̭EQ��n4��y�ۤ�M�^t���s�	$�䌘��������ۖB�܅Y̻s�:�� ���S���$��ݔ�9��|�<R��Y0�������Y�}���!%�����������2��ν�m5j��٥$��,����s1��9���ٕ|m��d��Z�9�Y�z���%:[QD��3�҉>0�,)]�Su��h������<�8Lr���9��ym��@�^��x�8P��}ff��h?�?����o�Կ�w{ߚF&,F�Uqm��s����~JɆ@CP����)�ԏd��ź
��a?ǘ�DP��s��(�o|�:G>g&�k�C\�����n�U	E�dn�A;����0{�]ci��K�Y�;V`_mS
+7�<̟�t�n�VיZ�!�ƹ����=i;��Xv��ˑ�~hA�a��$���7y�O�e�n%�5�gk��E�Zs��F�hŴƄ	e���������.�lh����ܽ��\��d]+��2g��[G��)��R�\"�������X:��UŲj386tL���[VYl�!���Iz��ܕ�#�q�\�Nv�ġ�?�0�����v0S;��֐ۥ?k��9�*��Y݇('3�ja.J��ü��h��ӹ�{�/z�)X������!L�-��!�C(,�s{Y8qv����C��	ٿ|�)}
�9�9a���A�i������?��!��N�}1�0
��#=��4��i1���3$#����H���#ՕZ��u��o�z�0�n�����l�h�W�;V6f>7Z�'}���\}r�/e�Å#zQZҒ"��}��bI���w��-���ah�;�-eda1��B�!˞�X��i�"/���>�8ړN��G�D-af1/H�C8��h,.�n�	�]朇4a��;"�sY+��*���*-��,�#ŕi������H>OLyu�$�*����F�ʄ3�S���c�����B�"��{6��e���� P�yżY���(��������3����oCV�߈
Ψ�c:�"���=J���ފĊ���jLC���S�ق}����ԙ	�����F��pW���aPeg�޳�l�%A+��
j�����*��I0�F��x+O���F8�W���� ��+�Bf\n���ɲl��k}� Mv0�Ȕ�H58�Z��B��$tC�H.���j��s�W�au�NS�^��+ޕ�7i��?ri�{���A��B}�bRB�=AΥ���8���D��0v��αZߞ�.�,�kX1��ײ��ް�����E󉈎�'p��|�Q��`��A�4h�'�0w��+ƀ����{��<���os"?��<f ��G�~٫�$c��ރ�ԑ�q	8n��=�g��	V����Liɏ<,���:�,CFؕ<( �������O�(c�̰=]���E�`;�n(�N(7�>���'�$����WN�_�5
,��H��P�5䌙d��[U��I^Eh@��j��>��ڴz��ܹɶQ�����;,��k6�C�ۋ�T��~ׅ�k�{%t�׿��t~�6�������zv�=�%��j�."�y&:��#|-��|y���=�C��e�j=�7��8��.4�ۮ�x�q�����L7���4����D�J��$��[1+	�.=Nc�Le��w�:�kEܼ���a�
{����y�f��jmd%X��W�ׅy�̥�xH�})l��� �C�1ё�c��fH|�2JJ�F�G�?Y�:ɷ�d[��`����W�PR�Q�?z����]'"�O�H^�Ӥg;N���L��"*�-n����7�$��L��J�N�v@t���2_	~��"HZ;��l
���mo;t�儼;+����Rf�M;݇���GJ��BI�8IJ2Ze��T�xA�t��z�g�gi�����m��:R���_���97�u5���H��mS=E��.+���m>��K��,D��60��-zP���kLR�,�����4Z�Z�{��=�-W���DQh6��2�!��#� ��K1��e*�m��mu�zNǶ�,�@�u���Q(?��n�G$�9�g��(�Tr�h�5���<!��i8=�H,\<"����֚�5ZֈGIYi�J���<ۯ����Zm�y�kkf����rst��	�I�0d����z�bw�K�N��؁i?k"kE�\m����D�&
6�>���8�A��)����n�S,h�~D-�#�^�����X�؜I�6>S���r��0uQ�,3������[�jF�2��4�\Z΀���(���5	�]�$��@-!s�z:i}���7�����ʫ9"�R|��-򨩐�vT
K_�k�VO4c����X�oqV҈F�L$htu��`~���������c���N*��p��om�0a�މ���3�\�M��	��vH=Yh�p��A�6����,0{�$/�ș���ųNc���!��ZY蹻FȮ.I6&^�ç��V���<����Oz��a��[�q�F+��{k�B�=����[tS\tr�ᙎSO�N��q��K�V����h1��_����o\��4*|�S;p�PD2�_��'����y"��B�(=#��.��_ �>|N�ރ@{*g�5�H��iC��F�ء�a�R��c�X$.t�8�ծW(��t�E�7W���AO����&r�MYy$O�^������ʨ��ՓL�Q�)Ҵ�d*Ě�Ӗ�Q�tY�l��J��D��?'& ��=��ڀ�)J�b�u[�6������A���q�|t��^�)zV���o8=)��LنA7�j��pÔ�)�s-���Y���+޼5rʷ�T7��t���Ѱl�S>�
���Uf��io;�r�Ԩ{-ˆ���s�0����������RTh�ăa�٩C�bE*�}���X��c͙�z�P�T��ʞ�����;9�+d���<IG�a����NJ� ���9D�3YG����u�ֈs,_���O����nTn=��������	H�VO��+z��x�u2�����FUL4*$�l0j9{��f"փ��)�
�)��P�}���Z:8�6��t�O� ]�����߯�;�'&�7M��U�	��K��t�u�岟^�`�}9@£?�K,�5��Nх7v�GD�(󪹆͆��7<#�d����Z��ۤv�m������"M����q1Y�qJT;�F� �������\�k��zH�L�8Z*���+�c�ҁ�K���`�J��6ts締^�fh����gpc��l<�SH�`����%���B�t!�"��RAU�FZn�C�Ǐ�R����R ��1���G�<7�lQ������J8����\U��|-}ݽ���;�t��0�*��*_�5���4
��a ��ջ���O嬱Z��S����y�����w�c�u��}y1��IC�K�t��'�[�k�*9I�Z����<%P���Y iӟ��$y+����܋X��I�,���a������?�\~�d�~��L��3�d�>�p���ф���d�8q��h�I�'��\(�JQ�
���6[�(W��f���Y$��bX`a}s�a]�e��Fɺ)�@
���0-%R|rд�b����%���E@K}�?R�ٖ�G��@_��7�:���-9r��QF@���l���b��*�i�l#���8���	�hOiH�iX|q�/T�����PO�U�`B��ƴ%ք��M����D1	���=�v���7CA�X����T_��OV�I#΃<沽 ���� ���&J�s�/Д�o��/�ol�r�8�]�vt^v��GoE��ޒI��Z�۲�S^HJ�}�sW��}|�8�;�ՅB����d1&�������w�D]��:[ϭ,c�#M��ˣ^�Z�
���a�=6=o��S����5��)�^����xӊ��*n�~��H���\����Z@=���$���@7Pt#A��X6�sߥ�>P9~�E�܂wx�>�g&��x,x�ixT���\�On�|����M��͐�X���0վ�Ɖ���SFH,k<T�i��s���0��͍��O�}F��p
b��-�?<�࢞�)�P����QO�,B�M콣�M1֠Y����A��P�	V�
0O��c��ӈ��8��@9�q�|wW�3{6S`������f\v�u@;r���9���m�Pšq�첢��0��N��q-&��#3/3up��l)�lȾ�++Kg7�i�;Mӵ��T�h���	��������]��CG��j��:�	�16/�$@�+AI���ʀԚE�������v�}ڞO�ܠT�	�~~gK��+���XlxVHYEB    a482     f40|�r��q�?��.�#+0�!�LecˤS^��!�ƹ1"e�w_���Oe�9y>��^H#��4��u�b?@ҝ�Ȳ)	A���ye�jH<��s��t��ϝ�F���(�O[3���u�Ѯ���U��8� �ݡ�����ݗӹ��v����#���(�p�\@`_�n�B�J�Œ�����cN�Ȉ�y|m
$��I��o��8�},�k�����;ıC2�Z���A�Y z�}��A_��O������3��69�{��:9(��z���K�'Q�Kޘ�z W���)hW��כNo��:L�.��*s-#D#��~CՄ��%^b0�p�Q'��+�e�j�Ppk\�(p� @Q�`��Kڹ)b�#�W�1��|hڄ3����|��!@Q�T��]i�)��j� �/}���C
KL��py�k�5�����ę�Q�M҉M)%�`)k�lAXM�GE�Hl瑚�ߺ������}���5�Y���'�A��ؒ�^l�5cm�i��1�jA@čit�24����wX�t����	��w����ͯ��g����px.w�������M?�{�f}�s� >�		i1�	�R<[�\���|�Փ��GBlo<��_dOGn3o��0��E����m�3�V,�Z`C&[D��g�a���'q ѐ��~�]�τBxx�6�X�bE��� ��pk���S�cV�6��M�+��@�_2���±h�jx��x�9�J����L"�)N��X�1 +(~4���r����zÛP�#G�a�����?���!���Aa����@/3��W�m]I
���IÙ���������i�A'��B�om\ۓX�E�뭺ӽ��)&��,�s�KԞ0P�w�¬#M���KV0�/�
�r� ����q������DmPx�T.��[A��F�+�!Y�'ې��A4tvBV�l/$X��1��H�lj��!ŭZ�iH�
��|�giQY�mE;1ǑI�Go��U�R'r��f��h"�=.��6 �w�J�l����hq�P��G��2�(��cg%x�z��II�x��� ����=��\`-&���:Mr�7�U�Qc'����i���b5�7�ʘb��:�)������'�>t.2F��jy+���WL'e�?�_�f�����ٜ'���5��)�Wv���ZE�N��s{5�[35n��>>�)|[�z!��,�f�i
Ձ�V����Ws%�%J���v�R�4vM�����J7~e��	?�uy�+��\�E4n���ϕe�&�3��:Uq_�:�P�E��U>�A��rV�+�V���3'1��<���*��Q(9����=4~QR�Ss�����ߨ�ulZ�ˬ�x�+�c�ӭ�iГO��o��,Qe���O��	� �u{�K�BsSX�#k���e��ˏ#L��4 N=�M�TXH��g�l��o�\����>/j�����<ڰ/tm���KF�5��ߔV�Z�0h?���9���v͙�f�(�����KT�c2P��mgx��'��W��)�.���@��D9��¨�;�Aލ���T�Y�B�i"|:��27�DZ:Ϧ��I�����y���p8ě��^��~!�Z� �����&K����Dp�<���`�bK���*'$�a��1^h� I���R��F��n�v�~�'D���|�۫��Bl��%ǡ}�Jξ���-g��̳�_���A�eÓ��A��1$�2�=���גf��xIC���d��Z�J�8%Y9�*�g�g-�3��%�F�
=O�k�ӱ�S-�]�`��X#��(����H�����躐mEj�k�q��9�w�Q$R����!$�a�cGfڠ��,裢�rü9o���x��6]g�f��#����\*$�%9�R�7�O�V7�A]�}k���bL>��P��OS@�UՋiٳ0��ܷq��'� �5?$ό�$X������4�j2&m��p ��(P�X����^��&a��pj@�]�)���1*������:	���Q�w�U���֞�G^޽�����^�m��ǎ痺�r_#L	*���D��ټ���Ty��Q[wFo��S�H4]��މ�dZ�������1�� ҕ|��'��>��-%,�h�Mqco�$��?Ȭ�D�$��8h�d��L�'d���s ό�3�n��?�n��Y�x�_�$�-۔����WQ��I% �`���Q�(V|e���Ԙ�=s3IEgbE��F����Q��*r_���O��!�2 �㬎ٚ�w|�A�jֺX��#�'�ݕ_y^$}�Nk��Yh������Wݓ�@��&�#��+4��&�8�՜�Fu��S����q��U��GD��\`&13A��u�)t��ec�G��v�P\R�M�!�mx����z�D�1?5��QbjIZU�rƒ�����Jp.ZEV��1�;��P�n F�k�t�f?m��R�ۼc���Aa�b��-<7�3ŋ�����LQ}�s(���]�6�("�U�*��*�{��("���vB�k�V��v�T㳮����(\_ɩ�߭��M�l���'e���X��!ثt:���ǻ� ����{�t�|�X��*�=��Q��K �gJ��8}�1p��0�eiJ�5�NG�^�71�*��4Na��|LZ���C���*�%!�i��Iq�^ÿ��7Z҃^�#k�n?S��e��z�x Մ�$���r剪Fݨ�|����Z��Q�Ҡ{3��͌�X4�U`�������tE�B��@���r��6/��`^��O�7P�y�q-vX�P�;sψ(�N�K8��j75����E�l"��OwEr�ފ������%шA�]Z:�N���{������On�����3 ($@��,� d�,Ur?���#@B�5����$c�2f�R����C��J�	�a �TG���yh�!1�%�!A�g�����Q�Et�Z�q�Y�7��B3'�a>+�ME���~C�^ d>��|@�@�������V�BX)Է�jq�=��=YFʂ���.��䱡��+,���I��n%z~�<E�G�������[��]l�/׆J����"�Sj��q�N. ����~�u�s�Ɠ���jY�A�����
E�a��^ء�Hf��I�T 
B����n��X��p`���a-��%�$��/�����=��b�Y3�(B�>'�P��ʥJ�0����M�-����Y�&��� UnP �Vd��c�
u�Þ-x�D[c��u��v��� $S�c�0Pm�WVO��CS$i$W��r�"���.��v�R���=A#@`��5�O�j��ލ.�1Շ�$*�攓�/4�VL"j�ф��,Ret����V�:� �����X�y����[�d7���z��)�;��ԷW�U83�iL�M��u�H�sz�m��y�Y�.�J_F�B���i�U<kn_�\�D�I��+��E�p;w��ג�"�s�ʭ�ў���
t��}������]б#	S�*Aa��}�2�����_�dX�d�AY^y��d���h���`���o���iD
�d��}`�z]��K���Iz@z���po�H7%;�晚�\b�+Rm��|�"����r��p�=R����6jvb��SSXP0�`S��^��1�� P��ޱ�
X������,�^TYVp4:cESv�����|P߮���X=�o���o���5�C�QN�y� �ਜ਼��RҮ��u��F�]�3ˎ�e(��b�$���c����-J���W��_��xs�\7��Mi��\5_���n/�H��a2���﷝�IW�J!|?��_�T��J?�@I�1���%D!���y�:�Py|zG�?c2�ͺ]:_�z�8�?