XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%]�:�����l�ߵ���Jِ�����zZ��SʯSq�G�'�A��D#�H0�\�-c�C�J��n��@�I$N��O% EG����g~��mÐ��K�Z�k��	�`�I˯��O|{���tfϐ�6=�/{�c}E:� y��k-������b&I꠷s9��k��юk)���%�9��v�g(�jn�ϛ�q�3�|vT�yD��,��@-��3��Czt����l��n'�"~�cL�XA��3���\J0�j�v��a�io>�3�S�S�g{F��@Q�����Y�w�=κΪ��'l6�'X<*��m �ӕZ��K�� �+%�?M>/��DD�Ƹ�/���&����6r�����~���0'A6���8�:5��5,������:�/�����xa��;g��v��[D����&�]3�l�d���&Q�E$w�Y�x㎯$�p�𳨺&٘_M�_��Do���۱#�?�C���1�]�#XkP�>Y�xg������.��1�?�֟�����cK��U�& ��;�4��f\?�W���*�u��X�ȇX�?�6/�Bs�mb�d޻_mKn�F*	~�TN����a*�|3��q����D9Np�TO	�Ԡg76���#mT������q9�K1ӕ�0�"���Z�B�4�9�:�x���'�=��S�3� 3=��^N%�&<[0�غ����7����tZ��>�df�>z�:�?rRV3>:�ʲ������mfv9h�8&�XlxVHYEB    2639     7f0��0�W�"N9��џ���ј9b*�ǔ@��gN`��g�h�GǅW��mD�nql�?�>�ھ]�1��,���y*%!�L��?�)ި
JƗ�<�[�>9o:��0�s���{o�G��DL���ÿ�L���^�s�ry�}r`��MP#����Y�J����
L�8�:�o��#D�r�:�O�7���.��s�7J^'�H�E�� (h��[�0��V���A�Z�G�k.x5�9����9����jNٔ�3q��Z��������X�M�u�GO��;��q����0劽���w�4-nţɄ���%և�tb��*m@sw��$�V�؞�d��*z�������� X�a�}���F���=d�fƮ ���M���v%<��ه��'晗���%kd<�<0]���]���/0ٷJ�C{Y�{Z)�(�R<��=,��B�FIyI�t�L�V�s��y�����ƪx^����./�4"iz~��=
�n�_i�P�Jr������N�g��#wef��)��Ug[%�k�������K�c#�`�lv+�G�;��}����� i��?c8_+3�/�o�=��5o<m�e5I,�!Oy�SZZF���fr�e�:Mj:Kg�����\=u'(+���@��F�V��Б�5�dǩO���M�/�V��ҍ|�\F91i�f%V��G�ۦ2�|��N\��$�l��\�	�];��_S�І��?.�hT��<3G��kPΜ{������vz׮�ϣ���-�P�\&Һ��_,��S �K���Q;�G���ߜ�o\��\� �{ā"7�)�ǝ��g����(�H��j���f�[��Z&	N��9Oa�q:�9�?�L��.��,4�{������%�#u:��[�@a��T�]���
.4C��N��3�@��b��#3_�0(�.˶������q׿t��>A�c�*�G*+���r9Ѻ�<sD���������� Bʡl��V��D��a�}��֖�n���/�1Μ�c�8�^��W��G,X��2ڑi\��Al��Ǥ�;��|Y�d�y�g����K�3l�����d����=҇A�0�0&�����.��m���Ha�%ߋ���^@���@c�!Y�M�x??,Ft��:�݇��#�v�Zl=����7<6�����%�� �^�6��ySF��sT�L\�:���G�*49�j+�JY�5�:��w�H~`�b9/��.�²$��Sb[�50��?�/[V���ʔ��2[.�v�J�N�c&�����@�m�h���.w:dKSU��Loc:;���m1'!5�@��OϮILr_Z���M�T��Q���A� ?�<~�RmlU� ݧ�^��[��sX	�2�n�QN��2�;L��2.&���np*Tع&@n$��e��;�4.��>I���Ia`��P���,�s����g�=���5P|^�`3�����ۓ?��p����z��d<�s �F��/<qG�>�����E(�9Đ��Ί�[la�@;�v�I�oR�>���~�Ps~�*�^��cv�c�<��;�HW��e	􎊫�ĉ�]/��|s�t^�ھ��T��摨����L�5�KCRMxw�S ��hZC	�&��J�\f�o��E�rG��m��fu���-!�~d�s�ה�0j��Ё�;D����\��`�Dkm�B�WS�j/z��o�Z��*Z�5p�I�+���K��K��V��x�%�kJ�@�a�$���I��oq�ה�L4��1ς��M�����+ �/׹H�CjΗu4`����qp�@����N��W��E���K�-t�m���K��G�ODE����`(#�JwӦ��*2��L��0a��Nvj����HR�E;M���l�b��]�6��cuz��摔�N�D�s��'�[癩H���4�6��O��>�S�����=��2O�@��G����.;���iL��>Tc֛���Ʉ��t�	�X!�����#��~�