XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������Y�����;����	O��"p+Ix]��I@J�Y�isy�ܷ �w�vF�Yu�Ӂ&F'�Lj"S4fc���"�5;��j�7�Ke����t��!ג�3��Ɠq0x,,x��&�iI0>q'M!`��󇨪��ۺ�>8�� �)I
����xi!�a)�1�u|6l�Ŭ�s9���k�,G,��s;�ΌL�E��t�:�qX���\C�4�����������ǖP�Ԅ�""Y�{��$��uV���Ȳ�:Q5.�9������� ��3s4fB㙆�i��y\H��x<])C���\L�5:�k�@f�9׍>��Ҩn�+�I���5��x�gX�;�o�ɞ�GI�W��_R��<2t��.6����񸇚Dl/	����0a��.9��&NE�R�Rm4���O��{���Q&ω)�=%��H�K��̽`T�@3�xس1�z�9f��(��4���s�u����L�Kr�b�C�?N��
�$�2҅����z���a��r�1����Im���J;�i��Q��0j��K˧��Y�%�>�V�y��R� gg�é���k�f�J����/ej�ío�n1��q�e�e2�x��ł���W���L���FfED��p-BgZ��pL�j�8����$vꚥ� fy$�!��oݾ�44=����v^���ig�*ęB�%˗��~�L	}τ������>�T�(f��� ��\j�>��ud������}*�hI؋�d�fK���A�<7'XlxVHYEB    2c4c     7a0�A�J����\Dn��R!��{�C��i
�1Q��|;n�!���O��Bk�R�W��m�8�N!G��o� ����5���,3��������c��<�-Nt�� �N4Y���#瀄�������j6jРV���?'�K+KJ�f�$o���J=I$b;��ǿ���Ӭ���"������^�KW'�T���yr��:6:_�@x��}+)�AEP�#�X�E��t�x��BB7��P����oO�u�n�bZ�8���V��R��_st<X�8��^&Sf<P�C�)��B�6���݉��u]/�;��B�şB[�P/�W1y`-��wI����l�0�,,Kc�`-<��=��EϢO٢y��"Ǝ�I2"�s���`���щ��������v���	-�m��9Ոt2Bs��[]�5�G���d�؉�}6B�S#�W;��V�J�| WᖁÒo����$QZ}J� G��D�vd��ҩz�L�z<{�e�|�c9��22?ﻦ�xj!�_�$�3�ޮ��=�7z�A�����{l�||��� ~�W����'f
7�,��h�޷Snct��Ȑ4��ӣEZױ�PfZ��x��Wc�f�f�^Q|ѤP@����F���!4{�Rzb.���g�(�QU*c�ZEk�	��Ǳm�D�""�n->D�m�p����y�x�X8��(��j���}ø�����<$��P��KVsy�B,�%��߄�m�P^��M��S"O��B�z�W��2�`�>���xI.�&[Ƕچl�7L��;0�ż�x񒜪	��������(E��~��n�<P���R���}��+Qr��Y
���4�m�
uf�NSc���}R��v��%��ZOWE2�-�-]l�vO�B�i�p&fD̸<���䅠�)�����|8Ҋ���p�'{#�%P_�ťЧ�b��E��� ��n���[��XxT1���y�f�؆����L��c*" ��c,tmK44-��(W�4��к�= P�*�%�y��ʆ%P�(B
��1:��较�Φ�0���_j⒧.�k����Tu�_3tS�VF��ݤ"�# `�~���.'Cq�B�I���
�(!u�U�B��f����!�?S����p��������ގ�y�wc!���rs���ۆ�֚����>c
E��ca�jJQ�'������J$���7��a*��dy���fë�I���~
e,	5z��=�R>�!LS���'���i��b<N����&��kG���jo�t�ӾAq�AY/Xx��0yn- 1p:0�� ����2jOo�]�mjrTVō0�x���卻���X�X���%<oڪ����	[�us��7�`G$yn�U+/�Á�N����Q0�(�k�*"�#�o�;�h'̻��q'rW���s&������ 	�`��@�4�S\SnN܏0x:ˈln�S���C_�-�ӌ��C��	P�O��,�;�4�i���P� I.���;�lHn���0�X̭����c�'0��}z��̕����өe�Q[5�FY��0[�ε�,�%ت��l��M��o�c��K��?bA�CK3|7B���%��Y�kz=��2�=ݷ�qR�髀2�vw��BIY�*(����I��b�9%��Q�ʼ�$��a���2r�_��0�}V�?�ڤ/�7)m���F]��t�K	.��/R�����-�q�D`�*���$��K���5���:�@H�B�9[�'o9P��f��Y$�rt�l�0g���@��]9=`"�Nvsc+_�����1��a��4nB��:���R00>4l�/��WG�`�F$|֮)�=��%��<Rt���;�C]чA|G���/Y���ZJ	ɮvZ�>����tU��Ar@{.��#��8M�>�?Ԅ��S���q��S�щ�|���]��dZe��K