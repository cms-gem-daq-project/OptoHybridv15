XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M$2��-�IQ���?߭`yݣ�GDw[zPG� u2vk
5��R��'se7w��5n`芗�������Lb<�%l��+5��k���n~êo�y��\����9�f]d-�@�Xb�䟈��ItN}�#�s��)��C7�4'y��k�iï$� �XW�T4�q��P�p.��p��ҤGΰ��|���zSFKx�%��M�K6*�;:�g�9��`0E�󮊯�V�.'�}7�+�<֡��x�G;�^NH\4�!�qޤ, �}qqs���ʶ��e�$'���Od�Ѽ����b�~�E��'�/f�q*94+�����3�i��^�o�Z��:��j.fJ���/m�O��i�cVCW���(�n�.�g��i�dJ���j����N�����oL	F%�<U!z��Q��L�� � �(�~:��mx�1޷�����CE�+�L���Ɋ�!GC���V�;���"�>��90�z�V�NI��11�����h��U�`/����� ��4!h�O�3��A�TO����L=�V�\=6�)K����N���������5��FE��kG�˴���rC�^�i;iX�K�P���eWN�d�)�.��]�ѱk�N%��5.6~gF�i�@�8Z�y.B	2����%%-���W�dUb#���䂰S����8Օ���T����@F������VL<z&��rt/]rE:�z�Pf�}��Kݸ��89�&�_���[&#<�b�m>��8�����%��^�FO4�q�XlxVHYEB    17a1     680�_ڂ�`\�r/^|��Ǌ�@�A3W��W����>�/�	�/��&��K t�q}e���&5N���W��tw
�8��;���>*���S@���R��^pp4�^"NC�@�Dq}�����H(A�N�Tr�~��枈��ԣ�]v*#./Q�R�͖��@[��[�M�羊E�&�R�F�ާ%v�	��v���N�C�Ϯ�qσ��8A��l'��dK�~���]D��lS��q��3kX��4=H��Z(��U�mdqs xY�uC�
A6S��gnڸ�~@��	[�N��r�=�~�N�`F\�d[�
a�rEC��!*0,��L�k�w��>hYal�};'m��)X4�m/�p�钮��ߗ�Pc��E�|��)"�,��<�D{�h�5���r���t�w�ڏ���j@De��Γ�9�C'ǈS[|
��K9c�-W"�BfU�Cs���X�E�n��t�银�� �[i�����Ps���$�����E�
�sZK������a��w4ġPΆ�}A	��6�c�10�`Sw�j�&��keyP���-8���jc���Ȕ6��¸�Ukհ��s�il��@�� �go5[���	�ӐAԶuj�*��Z>��Qg��/��M���r�H�k�J��I�g�0�*l?����6K�?5]���+Ց�Ӌ�����$��K�-+b���<��sm��6���)(8w!�R x��<?����	25_���B������nߔ I�b�Xg�𱩲�&��P�ݎ����2`��i٫T�;o��V��#�y�ɦt�rX��9`h�����kC�
� J�]�4i=��&��?K�J>�k?�*(�	x�:�T�sW���P)r���E�/�������ƑT����8⎎m��/~�"i�w#.T�7�hިX]��)8M�߶8'+툻c�~�1��9� 15�J�4��B^E��_6T�,4*'�V�Jb�&�K�]]n/��d���(q�������l��^�m<��>#m]iP��!�1_;����8�./��g�\���iFg�-�RF@|������jx:i�"r�׆���Y�n3,����+�C�}'��B`c����6�xd���2� ^>����+C8����\�����i��d\]�NdAyC*���G!YTn�C������Wzx�3�}��?���DK�]�Sj���U�b�2e'w�r��_R�T������EF�\���'�X��5}��w��(����ɾX� �\�2G��S��( A�� T�<�����H�������7�Pg��95B�����,I�,�Wm�X;���@z1�N�'G�6h���+d!5��u�Ԭ��!�`Y陸�����S R�jvP}�$i|{����}�Z1��4��fp�Kwo�?�'��^��/Y�$�8�O� 	���$,�6b�"�"�3*c0���s�10�&'�,��������8=0�\�-�����8��|�(�oLR�v��E�`������2TRW�$)J���a�4���梎����BԌ��L������<}��3^|LD��}�����
���wL3����o�g����ŰⲢ�dR�Y?�����m��g��4���J���
�����n�JnR�8�/d�H��