XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����U��=/�@�WT"Cv�뇓[��S���u�X��f��f�9o�m� 5>�0�O������"�
ݼ��*�;�Р/E��~v��[����P	>-�N��ϓ���H(�o�qu�N�H�]97;[�np�`R��0��~z[�ۚ'V�Ό��U9Cɞ����c'��x?U�q<p�&�|�Om��57�)Q�e��gj���ێ�~(��ca�b�%L'G]1&����ڏ*Q���!$�s�T�� S�_�1����q�\�-��W�U�M�����{4�5�=\�y S^l3nG�)dq�R�	��_��k���X����=1Bt���3L�$r�{&1a��خ��qr2�����߬!�4���0�g�#����wNX�����R�I���*f7�2��H���>x��^qbW�(�qO���B	��tp������x����|�Wy��`?�@M 8	Z���e�Re3dޒ�i􍘣(-�o
���$�)L/.�;��$m�2����^`�ܼ��O6�h�M�q�ꮗ'O	��ȷ@����73͚��H����G�͍���GQ���}�`���e���bN���v�E�A�p�7�2M��|�|�r�j�Y�N�u����y�������d�A�>gU��G%#����+���b�~1ޘ���=۱��3�7�⠜�Ǻ�DB�^tr�1��P���[&�yXrC�_�	jOBr�ؔ��+U��fǌ��Yد8���#�%���+c"%XlxVHYEB     935     3e0�!{K��kj7�E�ϯ�
�x�O.dX�,����@��e6����~*�ZX�Ƙ�z�YX`z��K���m�����9�$ X��p$}&�v<|�k��b��&lj[	��bh[k 1X<��@�)y�?z�1�NRW��q̂���A��l���%��XY�LQ��_�.,���5�� ��43�#���P�=u��	�N_
�����l���ָ�T~:�����EB�tf:���6f&�#*���ˇI�%��h��"O��^�h"9��3X��-�����	Ufu�4D�C�Y5rB��y�ؐ����a������=����2VqբyHB������9�t�1%ܛP��U��B$� o:��G>K�X��z�${U��gr�9w����D��Ψ�$/~#���@�7�zj�4�r������m��)��8��H�xx"�$��9{���	���	1+�o�6I&��H<�k���$��֌���v��絟C���ZN�
�bbpeŶUx(07 Km/�6��R�C�����bw	���Ҡ�U�dg�!����/�ؕd���GT�D�c(��'#�S�Sz������#ꢭ$��"�Y6�7L��܌�)M޻�pU�L�m㗡��ޜ���Uu���|�b4���c�Fi&���[���Q�z�sM���g����%�12����� �Bww3����{Q�U�3Tr��^��G�gV�1� [[�
?�ͼ�k����ko�ŤĂ0�tOwz��T'��_�� 8yx���6�]��L���!KHF������8P��4t��Z?ԅ@7�D�~F�a��S���էDT+3+F>���Uȃ��	R7* ����9Ձ2�x���!(|AA�����F�7�U�{��=��p�k�ׇ��4&f'��%�3�֠*9�Y;3}� �T������اґ�ZE(�p�?v��4��zd�N@��RV���^݈wؗyK����