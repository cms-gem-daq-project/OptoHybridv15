XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e�/��5���D1�PG�	r�,��7���P��� !ş��P�t�s��p̐e)�b�H�M1)�N��/��G�=n&��5��1�(M��C��t�]5�l��%� ,�y�G+���^CZ�>�m�o: ���)d?���<�!2�mڄ]��j�4��3
��FK��y�VŽR�����X����)h1�&nfG�t�~LׇR���[�/�$�b}���i��ڕ#�o�R��r�&�{�{`M^����-Eq�*ג}�<���a���L	�B��mƞ�@;�X�-҂�<X�H�#-L��܁H�@(�����dEc�<7%t���`�\�x����lhز=i-6j
T].�S�C��⻋�{&�[��)�a�3
%��d��8�Ү�����b���ĩ��$�̣��A��r�|K�Vu��
g�'`�)��
n"˼�Z6���Y����@��>k�P&]�a��X����9?kZf���0�X���Z��X��PF���-Kr`�DR�Q�$:���e��b���>���l�+�ѹntͪþe88, �0�n(���N�_������ߦ�㜉��Y��1͐4Ľm�xP�<�a��M��,B�L�=�)�Y�u��a�U�'࿜o����g����j��h\�$����U��r�f�/�v��<a$�"��yHRBϖ�rc^+p��n��w�s��(�֊�Wj��QY�<��m���׌=ei"�u�#�˒b��gD8�x.�b���H��"#y�d���^'��kᥦ�DXlxVHYEB    1cf8     790�t�!f
1O��~��ϡW�����|ģb>�m��@q�ɥ�z���o�q'Fm_쑂I���d1;a�������G�f�J���2���D����z��Äj�K��j_d�°//�������: �W�>�ƹ�r�]'h��u:���߷gs5+�q��ÀjF���8�37s�]��4�r��g�d�?��8_H�/���07}v$��ܟԉ@]vZn_*�1�7�%��p��W��4��ا�1� Z�h7�,�аp��!����r*Q�l:�" ���/�f�-�m
�;^�w�q�I{s����������lSFct]��"wϰW���vJ�S��/�=W��v��꽾q�`�ܕ�WV�[�`�ɎmQɌc^�u���߃�p��oe�^/��:�k[UrFR� �Rl��e+���L;� ?�H�T=�5����ݑߩ<�qքA�Q�S��CL�L/u�����E6����h>Lr�s�3s�ZA�r�Ne��ǥ4G8du:~�-�֌�@֓t�����e��X>��t���§
�[���G���v�X�s��&�۲2�"�}������3�����m��\�ӧS%�"�ʒ/��Q��<ODbt%��6�-m���;�A�~4h2T���y'jfcO#~Y�V�,���R�:������ɰ�%ǜm��*a1N�������,�4������x���e��SM�Cu�`��}��o��M+�%��a��ζ 8�omޮ1��/!�:���2�j������6q��kIt�A�:ΟZ(��Mw�c�2������0��QrByb���l��U�5t���i��@�w�Zf�`��h'k�AF�5������ᚣ�b���Lѓ=}FD�L�g�^�;"������T��G���1�f�SX��K���s��7�"kGG��a,ڰ��'=5I9
k�`�[������J$?�@���n�!��XeD�$*�G�_=!6�9" �S�v�?���5�k��E���A�}oz%�nݷ����E^7�rP��'N$��s�"%k�N؆�Q7�6q�*9���-Jx���:;[,����r�A�<����2�{~�|
���_�\�s�-��׺����mb��tP�������������Dɬ��>N=RZB����>M��9��@��m鑐F�Ň�TO�E��p�zn�እ3��)MJ�}Z���B68m��\�־҃P�N�b`�.���f
gL���:��pK����S� �y��{+=9��â����m�y��OC���5����Z}Q��A�~�����8��hߒ���gܞT�	�)K5CТ}�x�O���!��W	ۻ1?�o(�w��F��؞�4a�5����2W�X�Ue<u���]2��Dߘ=��pW��@ڞ����mT��8����p�Em��X��	c�=�i������@���}y��f��@��l�]񇿷b�������b�Av挍r)�W�˒�Gz�c��85��_$o�w!�w� )��.�9+.����z�u�����|5����T�3�9<+Y9Eb��M�%V<r�j:��Z:x�l�F[�w������Dco���H�	 e�_�lzl(b�x�>d���J)��e*�`��<�@k8t���嚅P;�7]�:k$��_=�N�k9��OVT�S�g��EF7�����iH�,���0 ~M�d��g�=
{�b�h���syzÁɜ�_2��[��r�	�g����#�ϥ/�h�;S�[��!X�N�HZ�s��z;{;�x�V�P�IW�ޫ�T���ϤBN���/��Ip�t����у�*q��
����Yf�L|�J�0�$�E����Urs	v�C�l��5N�E�M���g,�l짠��.��$���&r`<